magic
tech c035u
timestamp 1386015194
<< nwell >>
rect 0 402 720 746
<< polysilicon >>
rect 216 681 221 697
rect 351 691 358 719
rect 381 691 388 719
rect 432 704 499 711
rect 28 671 35 679
rect 58 671 65 679
rect 88 671 95 679
rect 132 671 139 679
rect 162 671 169 679
rect 189 671 196 679
rect 216 671 223 681
rect 28 375 35 623
rect 58 553 65 623
rect 88 539 95 623
rect 132 553 139 623
rect 88 523 93 539
rect 58 381 65 505
rect 28 235 35 359
rect 58 335 65 365
rect 88 335 95 523
rect 132 381 139 505
rect 162 381 169 623
rect 189 501 196 623
rect 132 335 139 365
rect 88 319 93 335
rect 58 235 65 305
rect 88 235 95 319
rect 132 235 139 305
rect 162 235 169 365
rect 189 355 196 485
rect 189 235 196 339
rect 216 235 223 623
rect 318 610 325 621
rect 246 583 251 599
rect 246 553 253 583
rect 246 358 253 505
rect 318 388 325 562
rect 351 486 358 643
rect 381 612 388 643
rect 434 612 441 623
rect 475 612 482 645
rect 492 624 499 704
rect 537 691 544 719
rect 595 691 602 719
rect 537 624 544 643
rect 492 617 544 624
rect 537 612 544 617
rect 381 486 388 564
rect 434 486 441 564
rect 475 486 482 564
rect 537 486 544 564
rect 595 532 602 643
rect 663 612 670 675
rect 246 275 253 328
rect 251 259 253 275
rect 318 220 325 372
rect 351 331 358 438
rect 381 402 388 438
rect 434 428 441 438
rect 450 412 462 419
rect 381 395 422 402
rect 415 358 422 395
rect 455 358 462 412
rect 475 410 482 438
rect 537 428 544 438
rect 475 403 503 410
rect 496 358 503 403
rect 537 358 544 412
rect 351 288 358 315
rect 415 288 422 328
rect 28 197 35 205
rect 58 197 65 205
rect 88 197 95 205
rect 132 197 139 205
rect 162 197 169 205
rect 189 197 196 205
rect 216 197 223 205
rect 318 182 325 190
rect 351 161 358 258
rect 415 220 422 258
rect 455 220 462 328
rect 496 220 503 328
rect 537 255 544 328
rect 537 248 551 255
rect 537 225 551 232
rect 537 220 544 225
rect 595 220 602 516
rect 627 486 634 539
rect 627 358 634 438
rect 627 288 634 328
rect 351 110 358 131
rect 415 127 422 190
rect 455 128 462 190
rect 496 161 503 190
rect 537 161 544 190
rect 595 180 602 190
rect 595 142 602 150
rect 627 142 634 258
rect 663 227 670 564
rect 653 220 670 227
rect 660 190 667 195
rect 653 188 667 190
rect 660 180 667 188
rect 660 142 667 150
rect 496 120 503 131
rect 537 120 544 131
<< ndiffusion >>
rect 56 305 58 335
rect 65 305 67 335
rect 130 305 132 335
rect 139 305 141 335
rect 244 328 246 358
rect 253 328 255 358
rect 26 205 28 235
rect 35 205 58 235
rect 65 205 67 235
rect 83 205 88 235
rect 95 205 114 235
rect 130 205 132 235
rect 139 205 162 235
rect 169 205 171 235
rect 187 205 189 235
rect 196 205 216 235
rect 223 205 225 235
rect 410 328 415 358
rect 422 328 455 358
rect 462 328 469 358
rect 485 328 496 358
rect 503 328 537 358
rect 544 328 549 358
rect 346 258 351 288
rect 358 258 415 288
rect 422 258 433 288
rect 316 190 318 220
rect 325 190 330 220
rect 625 258 627 288
rect 634 258 640 288
rect 413 190 415 220
rect 422 190 455 220
rect 462 190 465 220
rect 529 190 537 220
rect 544 190 595 220
rect 602 190 606 220
rect 346 131 351 161
rect 358 131 363 161
rect 494 131 496 161
rect 503 131 537 161
rect 544 131 548 161
rect 657 150 660 180
rect 667 150 670 180
<< pdiffusion >>
rect 26 623 28 671
rect 35 623 40 671
rect 56 623 58 671
rect 65 623 67 671
rect 83 623 88 671
rect 95 623 114 671
rect 130 623 132 671
rect 139 623 141 671
rect 157 623 162 671
rect 169 623 171 671
rect 187 623 189 671
rect 196 623 198 671
rect 214 623 216 671
rect 223 623 225 671
rect 349 643 351 691
rect 358 643 360 691
rect 376 643 381 691
rect 388 643 390 691
rect 56 505 58 553
rect 65 505 67 553
rect 130 505 132 553
rect 139 505 141 553
rect 315 562 318 610
rect 325 562 330 610
rect 244 505 246 553
rect 253 505 255 553
rect 520 643 537 691
rect 544 643 554 691
rect 570 643 595 691
rect 602 643 605 691
rect 379 564 381 612
rect 388 564 416 612
rect 432 564 434 612
rect 441 564 451 612
rect 467 564 475 612
rect 482 564 484 612
rect 500 564 537 612
rect 544 564 546 612
rect 660 564 663 612
rect 670 564 680 612
rect 349 438 351 486
rect 358 438 361 486
rect 377 438 381 486
rect 388 438 390 486
rect 410 438 434 486
rect 441 438 449 486
rect 467 438 475 486
rect 482 438 484 486
rect 500 438 537 486
rect 544 438 547 486
rect 624 438 627 486
rect 634 438 640 486
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 174 86
rect 190 79 202 86
rect 218 79 230 86
rect 246 79 258 86
rect 274 79 294 86
rect 0 76 294 79
rect 310 76 322 86
rect 338 76 350 86
rect 366 76 378 86
rect 394 76 406 86
rect 422 76 434 86
rect 450 76 462 86
rect 478 76 490 86
rect 506 76 518 86
rect 535 76 547 86
rect 563 76 575 86
rect 591 76 603 86
rect 619 76 631 86
rect 648 76 660 86
rect 677 76 689 86
rect 706 76 720 86
<< nohmic >>
rect 0 743 294 746
rect 0 736 6 743
rect 22 736 34 743
rect 50 736 62 743
rect 78 736 90 743
rect 106 736 118 743
rect 134 736 146 743
rect 162 736 174 743
rect 190 736 202 743
rect 218 736 230 743
rect 246 736 258 743
rect 274 736 294 743
rect 310 736 322 746
rect 338 736 350 746
rect 366 736 378 746
rect 394 736 406 746
rect 422 736 434 746
rect 450 736 462 746
rect 478 736 490 746
rect 506 736 518 746
rect 534 736 546 746
rect 562 736 574 746
rect 590 736 602 746
rect 618 736 630 746
rect 646 736 658 746
rect 674 736 686 746
rect 702 736 720 746
<< ntransistor >>
rect 58 305 65 335
rect 132 305 139 335
rect 246 328 253 358
rect 28 205 35 235
rect 58 205 65 235
rect 88 205 95 235
rect 132 205 139 235
rect 162 205 169 235
rect 189 205 196 235
rect 216 205 223 235
rect 415 328 422 358
rect 455 328 462 358
rect 496 328 503 358
rect 537 328 544 358
rect 351 258 358 288
rect 415 258 422 288
rect 318 190 325 220
rect 627 258 634 288
rect 415 190 422 220
rect 455 190 462 220
rect 537 190 544 220
rect 595 190 602 220
rect 351 131 358 161
rect 496 131 503 161
rect 537 131 544 161
rect 660 150 667 180
<< ptransistor >>
rect 28 623 35 671
rect 58 623 65 671
rect 88 623 95 671
rect 132 623 139 671
rect 162 623 169 671
rect 189 623 196 671
rect 216 623 223 671
rect 351 643 358 691
rect 381 643 388 691
rect 58 505 65 553
rect 132 505 139 553
rect 318 562 325 610
rect 246 505 253 553
rect 537 643 544 691
rect 595 643 602 691
rect 381 564 388 612
rect 434 564 441 612
rect 475 564 482 612
rect 537 564 544 612
rect 663 564 670 612
rect 351 438 358 486
rect 381 438 388 486
rect 434 438 441 486
rect 475 438 482 486
rect 537 438 544 486
rect 627 438 634 486
<< polycontact >>
rect 221 681 237 697
rect 416 695 432 711
rect 466 645 482 661
rect 93 523 109 539
rect 24 359 40 375
rect 54 365 70 381
rect 180 485 196 501
rect 127 365 143 381
rect 158 365 174 381
rect 93 319 109 335
rect 180 339 196 355
rect 251 583 267 599
rect 654 675 670 691
rect 618 539 634 555
rect 590 516 606 532
rect 309 372 325 388
rect 235 259 251 275
rect 434 412 450 428
rect 537 412 553 428
rect 347 315 363 331
rect 539 232 555 248
rect 618 328 634 358
rect 487 190 503 220
rect 595 150 611 180
rect 644 190 660 220
rect 410 111 426 127
rect 451 111 468 128
<< ndiffcontact >>
rect 40 305 56 335
rect 67 305 83 335
rect 114 305 130 335
rect 141 305 157 335
rect 228 328 244 358
rect 255 328 271 358
rect 10 205 26 235
rect 67 205 83 235
rect 114 205 130 235
rect 171 205 187 235
rect 225 205 241 235
rect 394 328 410 358
rect 469 328 485 358
rect 549 328 565 358
rect 330 258 346 288
rect 433 258 449 288
rect 300 190 316 220
rect 330 190 346 220
rect 609 258 625 288
rect 640 258 656 288
rect 397 190 413 220
rect 465 190 481 220
rect 513 190 529 220
rect 606 190 622 220
rect 330 131 346 161
rect 363 131 379 161
rect 478 131 494 161
rect 548 131 564 161
rect 641 150 657 180
rect 670 150 686 180
<< pdiffcontact >>
rect 9 623 26 671
rect 40 623 56 671
rect 67 623 83 671
rect 114 623 130 671
rect 141 623 157 671
rect 171 623 187 671
rect 198 623 214 671
rect 225 623 241 671
rect 333 643 349 691
rect 360 643 376 691
rect 390 643 406 691
rect 40 505 56 553
rect 67 505 83 553
rect 114 505 130 553
rect 141 505 157 553
rect 299 562 315 610
rect 330 562 346 610
rect 228 505 244 553
rect 255 505 271 553
rect 504 643 520 691
rect 554 643 570 691
rect 605 643 621 691
rect 363 564 379 612
rect 416 564 432 612
rect 451 564 467 612
rect 484 564 500 612
rect 546 564 562 612
rect 644 564 660 612
rect 680 564 696 612
rect 333 438 349 486
rect 361 438 377 486
rect 390 438 410 486
rect 449 438 467 486
rect 484 438 500 486
rect 547 438 563 486
rect 608 438 624 486
rect 640 438 657 486
<< psubstratetap >>
rect 6 79 22 96
rect 34 79 50 96
rect 62 79 78 96
rect 90 79 106 96
rect 118 79 134 96
rect 146 79 162 96
rect 174 79 190 96
rect 202 79 218 96
rect 230 79 246 96
rect 258 79 274 96
rect 294 76 310 92
rect 322 76 338 92
rect 350 76 366 92
rect 378 76 394 92
rect 406 76 422 92
rect 434 76 450 92
rect 462 76 478 92
rect 490 76 506 92
rect 518 76 535 92
rect 547 76 563 92
rect 575 76 591 92
rect 603 76 619 92
rect 631 76 648 92
rect 660 76 677 92
rect 689 76 706 92
<< nsubstratetap >>
rect 6 727 22 743
rect 34 727 50 743
rect 62 727 78 743
rect 90 727 106 743
rect 118 727 134 743
rect 146 727 162 743
rect 174 727 190 743
rect 202 727 218 743
rect 230 727 246 743
rect 258 727 274 743
rect 294 730 310 746
rect 322 730 338 746
rect 350 730 366 746
rect 378 730 394 746
rect 406 730 422 746
rect 434 730 450 746
rect 462 730 478 746
rect 490 730 506 746
rect 518 730 534 746
rect 546 730 562 746
rect 574 730 590 746
rect 602 730 618 746
rect 630 730 646 746
rect 658 730 674 746
rect 686 730 702 746
<< metal1 >>
rect 0 782 720 792
rect 0 759 174 769
rect 252 759 598 769
rect 614 759 720 769
rect 0 743 294 746
rect 0 727 6 743
rect 22 727 34 743
rect 50 727 62 743
rect 78 727 90 743
rect 106 727 118 743
rect 134 727 146 743
rect 162 727 174 743
rect 190 727 202 743
rect 218 727 230 743
rect 246 727 258 743
rect 274 730 294 743
rect 310 730 322 746
rect 338 730 350 746
rect 366 730 378 746
rect 394 730 406 746
rect 422 730 434 746
rect 450 730 462 746
rect 478 730 490 746
rect 506 730 518 746
rect 534 730 546 746
rect 562 730 574 746
rect 590 730 602 746
rect 618 730 630 746
rect 646 730 658 746
rect 674 730 686 746
rect 702 730 720 746
rect 274 727 720 730
rect 0 721 720 727
rect 9 671 26 721
rect 67 671 83 721
rect 93 701 211 711
rect 15 573 26 623
rect 43 613 53 623
rect 93 613 103 701
rect 120 681 184 691
rect 120 671 130 681
rect 174 671 184 681
rect 201 671 211 701
rect 299 634 315 721
rect 333 691 349 721
rect 360 701 416 711
rect 360 691 376 701
rect 554 701 654 711
rect 554 691 570 701
rect 654 691 670 695
rect 299 633 316 634
rect 390 633 406 643
rect 43 603 103 613
rect 144 593 154 623
rect 174 613 184 623
rect 228 613 238 623
rect 174 603 238 613
rect 299 621 406 633
rect 416 645 466 655
rect 299 610 315 621
rect 363 612 379 621
rect 144 583 251 593
rect 15 563 238 573
rect 40 553 50 563
rect 145 553 157 563
rect 109 523 114 539
rect 228 553 238 563
rect 73 495 83 505
rect 73 485 180 495
rect 261 385 271 505
rect 299 511 315 562
rect 416 612 432 645
rect 504 633 520 643
rect 605 633 621 643
rect 680 633 696 721
rect 451 623 696 633
rect 451 612 467 623
rect 546 612 562 623
rect 680 612 696 623
rect 330 549 346 562
rect 416 549 432 564
rect 330 539 432 549
rect 484 554 500 564
rect 484 544 618 554
rect 390 516 550 526
rect 566 516 590 526
rect 644 526 660 564
rect 606 516 660 526
rect 299 501 377 511
rect 361 486 377 501
rect 390 486 410 516
rect 680 506 696 564
rect 449 496 563 506
rect 449 486 467 496
rect 547 486 563 496
rect 608 496 696 506
rect 608 486 624 496
rect 563 438 608 486
rect 333 428 349 438
rect 484 428 500 438
rect 640 428 657 438
rect 333 418 434 428
rect 450 418 500 428
rect 553 418 657 428
rect 348 390 485 402
rect 120 365 127 379
rect 261 375 309 385
rect 261 358 271 375
rect 73 345 180 355
rect 73 335 83 345
rect 109 319 114 335
rect 46 295 56 305
rect 147 295 157 305
rect 348 353 361 390
rect 469 358 485 390
rect 300 341 361 353
rect 228 295 238 328
rect 46 285 271 295
rect 13 265 235 275
rect 13 235 23 265
rect 70 245 150 255
rect 70 235 80 245
rect 114 101 130 205
rect 140 195 150 245
rect 174 235 184 265
rect 228 195 238 205
rect 140 185 238 195
rect 261 101 271 285
rect 300 288 316 341
rect 347 314 363 315
rect 565 328 618 358
rect 394 318 410 328
rect 394 308 686 318
rect 300 258 330 288
rect 449 278 609 288
rect 300 220 316 258
rect 330 247 346 258
rect 640 248 656 258
rect 330 235 529 247
rect 513 220 529 235
rect 555 232 656 248
rect 346 190 397 220
rect 481 190 487 220
rect 622 190 644 220
rect 300 161 316 190
rect 670 180 686 308
rect 300 131 330 161
rect 379 151 478 161
rect 611 150 641 180
rect 300 101 318 131
rect 409 111 410 127
rect 548 121 564 131
rect 468 111 564 121
rect 0 96 720 101
rect 0 79 6 96
rect 22 79 34 96
rect 50 79 62 96
rect 78 79 90 96
rect 106 79 118 96
rect 134 79 146 96
rect 162 79 174 96
rect 190 79 202 96
rect 218 79 230 96
rect 246 79 258 96
rect 274 92 720 96
rect 274 79 294 92
rect 0 76 294 79
rect 310 76 322 92
rect 338 76 350 92
rect 366 76 378 92
rect 394 76 406 92
rect 422 76 434 92
rect 450 76 462 92
rect 478 76 490 92
rect 506 76 518 92
rect 535 76 547 92
rect 563 76 575 92
rect 591 76 603 92
rect 619 76 631 92
rect 648 76 660 92
rect 677 76 689 92
rect 706 76 720 92
rect 0 53 347 63
rect 363 53 720 63
rect 0 30 106 40
rect 120 30 720 40
rect 0 7 393 17
rect 409 7 720 17
<< m2contact >>
rect 174 757 188 771
rect 238 758 252 772
rect 598 756 614 772
rect 237 683 251 697
rect 654 695 670 711
rect 550 516 566 532
rect 70 367 85 381
rect 106 365 120 379
rect 174 367 188 381
rect 24 345 38 359
rect 347 298 363 314
rect 393 111 409 127
rect 347 50 363 66
rect 106 28 120 42
rect 393 3 409 19
<< metal2 >>
rect 24 359 36 799
rect 72 381 84 799
rect 175 743 187 757
rect 174 727 187 743
rect 175 381 187 727
rect 239 697 251 758
rect 552 532 564 799
rect 600 772 612 799
rect 600 711 612 756
rect 600 695 654 711
rect 24 0 36 345
rect 72 0 84 367
rect 107 42 119 365
rect 347 66 363 298
rect 393 19 409 111
rect 552 0 564 516
rect 600 0 612 695
<< labels >>
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal2 24 799 36 799 5 D
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 53 0 63 3 Clock
rlabel metal2 24 0 36 0 1 D
rlabel metal2 72 0 84 0 1 Load
rlabel metal2 72 799 84 799 5 Load
rlabel metal2 552 799 564 799 5 nQ
rlabel metal2 552 0 564 0 1 nQ
rlabel metal2 600 799 612 799 5 Q
rlabel metal2 600 0 612 0 1 Q
rlabel metal1 720 782 720 792 7 ScanReturn
rlabel metal1 720 759 720 769 7 Q
rlabel metal1 720 76 720 101 7 GND!
rlabel metal1 720 53 720 63 7 Clock
rlabel metal1 720 30 720 40 7 Test
rlabel metal1 720 7 720 17 7 nReset
<< end >>
