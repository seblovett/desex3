magic
tech c035u
timestamp 1386006533
<< nwell >>
rect 0 402 133 746
<< polysilicon >>
rect 84 756 86 772
rect 79 480 86 756
rect 79 362 86 432
rect 79 324 86 332
<< ndiffusion >>
rect 77 332 79 362
rect 86 332 88 362
<< pdiffusion >>
rect 77 432 79 480
rect 86 432 88 480
<< pohmic >>
rect 0 76 54 86
rect 70 76 82 86
rect 98 76 120 86
<< nohmic >>
rect 0 736 58 746
rect 54 730 58 736
<< ntransistor >>
rect 79 332 86 362
<< ptransistor >>
rect 79 432 86 480
<< polycontact >>
rect 68 756 84 772
<< ndiffcontact >>
rect 61 332 77 362
rect 88 332 104 362
<< pdiffcontact >>
rect 61 432 77 480
rect 88 432 104 480
<< psubstratetap >>
rect 54 76 70 92
rect 82 76 98 92
<< nsubstratetap >>
rect 58 730 74 746
<< metal1 >>
rect 0 782 104 792
rect 0 759 68 769
rect 0 730 58 746
rect 74 730 77 746
rect 0 721 77 730
rect 61 480 77 721
rect 94 480 104 782
rect 94 362 104 432
rect 61 101 77 332
rect 0 92 120 101
rect 0 76 54 92
rect 70 76 82 92
rect 98 76 120 92
<< m2contact >>
rect 120 76 320 101
<< metal2 >>
rect 120 101 320 799
rect 120 0 320 76
<< labels >>
rlabel metal2 120 799 320 799 5 GND!
rlabel metal2 120 0 320 0 1 GND!
rlabel metal1 0 759 0 769 7 Scan
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 782 0 792 3 nScan
rlabel metal1 0 76 0 101 7 GND!
<< end >>
