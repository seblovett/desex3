magic
tech c035u
timestamp 1386266080
<< nwell >>
rect 0 401 480 799
<< pwell >>
rect 0 0 480 401
<< polysilicon >>
rect 183 538 190 546
rect 55 469 62 477
rect 153 469 160 477
rect 55 391 62 421
rect 153 404 160 421
rect 60 375 62 391
rect 55 340 62 375
rect 153 352 160 388
rect 183 378 190 490
rect 295 469 302 477
rect 415 469 422 477
rect 295 391 302 421
rect 415 391 422 421
rect 300 375 302 391
rect 420 375 422 391
rect 153 314 160 322
rect 55 302 62 310
rect 183 309 190 362
rect 295 340 302 375
rect 415 340 422 375
rect 295 302 302 310
rect 415 302 422 310
rect 183 271 190 279
<< ndiffusion >>
rect 53 310 55 340
rect 62 310 64 340
rect 151 322 153 352
rect 160 322 162 352
rect 293 310 295 340
rect 302 310 304 340
rect 413 310 415 340
rect 422 310 424 340
rect 181 279 183 309
rect 190 308 216 309
rect 190 279 200 308
<< pdiffusion >>
rect 178 490 183 538
rect 190 490 200 538
rect 53 421 55 469
rect 62 421 64 469
rect 151 421 153 469
rect 160 421 162 469
rect 293 421 295 469
rect 302 421 304 469
rect 413 421 415 469
rect 422 421 424 469
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 126 86
rect 142 76 154 86
rect 170 76 182 86
rect 198 76 210 86
rect 226 76 246 86
rect 262 76 274 86
rect 290 76 302 86
rect 318 76 330 86
rect 346 76 366 86
rect 382 76 394 86
rect 410 76 422 86
rect 438 76 450 86
rect 466 76 480 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
rect 50 736 62 746
rect 78 736 90 746
rect 106 736 126 746
rect 143 736 155 746
rect 172 736 184 746
rect 201 736 213 746
rect 230 736 246 746
rect 262 736 274 746
rect 290 736 302 746
rect 318 736 330 746
rect 346 736 366 746
rect 382 736 394 746
rect 410 736 422 746
rect 438 736 450 746
rect 466 736 480 746
<< ntransistor >>
rect 55 310 62 340
rect 153 322 160 352
rect 295 310 302 340
rect 415 310 422 340
rect 183 279 190 309
<< ptransistor >>
rect 183 490 190 538
rect 55 421 62 469
rect 153 421 160 469
rect 295 421 302 469
rect 415 421 422 469
<< polycontact >>
rect 44 375 60 391
rect 152 388 168 404
rect 174 362 190 378
rect 284 375 300 391
rect 404 375 420 391
<< ndiffcontact >>
rect 37 310 53 340
rect 64 310 80 340
rect 135 322 151 352
rect 162 322 178 352
rect 277 310 293 340
rect 304 310 320 340
rect 397 310 413 340
rect 424 310 440 340
rect 165 279 181 309
rect 200 279 216 308
<< pdiffcontact >>
rect 162 490 178 538
rect 200 490 216 538
rect 37 421 53 469
rect 64 421 80 469
rect 135 421 151 469
rect 162 421 178 469
rect 277 421 293 469
rect 304 421 320 469
rect 397 421 413 469
rect 424 421 440 469
<< psubstratetap >>
rect 37 281 53 297
rect 277 281 293 297
rect 397 281 413 297
rect 165 244 181 260
rect 165 216 181 232
rect 165 188 181 204
rect 165 160 181 176
rect 165 132 181 148
rect 165 104 181 120
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 126 76 142 92
rect 154 76 170 92
rect 182 76 198 92
rect 210 76 226 92
rect 246 76 262 92
rect 274 76 290 92
rect 302 76 318 92
rect 330 76 346 92
rect 366 76 382 92
rect 394 76 410 92
rect 422 76 438 92
rect 450 76 466 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
rect 62 730 78 746
rect 90 730 106 746
rect 126 730 143 746
rect 155 730 172 746
rect 184 730 201 746
rect 213 730 230 746
rect 246 730 262 746
rect 274 730 290 746
rect 302 730 318 746
rect 330 730 346 746
rect 366 730 382 746
rect 394 730 410 746
rect 422 730 438 746
rect 450 730 466 746
<< metal1 >>
rect 205 825 263 835
rect 277 825 383 835
rect 85 807 143 817
rect 0 782 480 792
rect 0 759 480 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 62 746
rect 78 730 90 746
rect 106 730 126 746
rect 143 730 155 746
rect 172 730 184 746
rect 201 730 213 746
rect 230 730 246 746
rect 262 730 274 746
rect 290 730 302 746
rect 318 730 330 746
rect 346 730 366 746
rect 382 730 394 746
rect 410 730 422 746
rect 438 730 450 746
rect 466 730 480 746
rect 0 721 480 730
rect 37 469 53 721
rect 162 538 178 721
rect 135 490 162 538
rect 135 469 151 490
rect 70 389 80 421
rect 178 378 188 469
rect 200 404 216 490
rect 277 469 293 721
rect 397 469 413 721
rect 70 340 80 375
rect 178 322 188 362
rect 37 297 53 310
rect 37 101 53 281
rect 135 309 151 322
rect 135 279 165 309
rect 200 308 216 388
rect 310 389 320 421
rect 430 389 440 421
rect 310 340 320 375
rect 430 340 440 375
rect 277 297 293 310
rect 165 260 181 279
rect 165 232 181 244
rect 165 204 181 216
rect 165 176 181 188
rect 165 148 181 160
rect 165 120 181 132
rect 165 101 181 104
rect 277 101 293 281
rect 397 297 413 310
rect 397 101 413 281
rect 0 92 480 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 126 92
rect 142 76 154 92
rect 170 76 182 92
rect 198 76 210 92
rect 226 76 246 92
rect 262 76 274 92
rect 290 76 302 92
rect 318 76 330 92
rect 346 76 366 92
rect 382 76 394 92
rect 410 76 422 92
rect 438 76 450 92
rect 466 76 480 92
rect 0 53 480 63
rect 0 30 480 40
rect 0 7 480 17
<< m2contact >>
rect 191 823 205 837
rect 263 823 277 837
rect 383 823 397 837
rect 70 806 85 820
rect 143 805 157 819
rect 30 376 44 390
rect 70 375 84 389
rect 136 388 152 404
rect 200 388 216 404
rect 270 376 284 390
rect 310 375 324 389
rect 390 376 404 390
rect 430 375 444 389
<< metal2 >>
rect 24 390 36 865
rect 144 819 156 865
rect 192 837 204 865
rect 24 376 30 390
rect 72 389 84 806
rect 144 404 156 805
rect 192 404 204 823
rect 24 0 36 376
rect 152 388 160 404
rect 192 388 200 404
rect 264 390 276 823
rect 72 0 84 375
rect 144 0 156 388
rect 192 0 204 388
rect 264 376 270 390
rect 312 389 324 799
rect 264 0 276 376
rect 312 0 324 375
rect 384 390 396 823
rect 384 376 390 390
rect 432 389 444 799
rect 384 0 396 376
rect 432 0 444 375
<< labels >>
rlabel metal1 480 721 480 746 7 Vdd!
rlabel metal1 480 759 480 769 7 Scan
rlabel metal1 480 782 480 792 6 ScanReturn
rlabel metal1 480 7 480 17 8 nReset
rlabel metal1 480 30 480 40 7 Test
rlabel metal1 480 53 480 63 7 Clock
rlabel metal1 480 76 480 101 7 GND!
rlabel metal2 24 865 36 865 5 nA
rlabel metal2 144 865 156 865 5 A
rlabel metal2 192 865 204 865 5 Y
<< end >>
