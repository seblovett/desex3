magic
tech c035u
timestamp 1386001875
<< nwell >>
rect 0 402 360 746
<< polysilicon >>
rect 44 672 49 685
rect 73 672 78 685
rect 44 631 51 672
rect 71 631 78 672
rect 91 631 98 695
rect 118 631 125 672
rect 148 631 155 670
rect 175 631 182 672
rect 206 631 213 695
rect 279 632 286 640
rect 44 504 51 583
rect 71 504 78 583
rect 91 504 98 583
rect 118 504 125 583
rect 44 261 51 456
rect 71 261 78 456
rect 91 261 98 456
rect 118 261 125 456
rect 148 287 155 583
rect 44 161 51 231
rect 71 161 78 231
rect 91 161 98 231
rect 118 161 125 231
rect 148 161 155 271
rect 175 161 182 583
rect 206 504 213 583
rect 279 550 286 584
rect 269 543 286 550
rect 206 261 213 456
rect 206 161 213 231
rect 262 207 269 537
rect 292 504 299 512
rect 292 287 299 456
rect 292 261 299 271
rect 292 223 299 231
rect 262 161 269 191
rect 44 123 51 131
rect 71 123 78 131
rect 91 123 98 131
rect 118 123 125 131
rect 148 123 155 131
rect 175 123 182 131
rect 206 123 213 131
rect 262 123 269 131
<< ndiffusion >>
rect 42 231 44 261
rect 51 231 53 261
rect 69 231 71 261
rect 78 231 91 261
rect 98 231 100 261
rect 116 231 118 261
rect 125 231 127 261
rect 204 231 206 261
rect 213 231 215 261
rect 290 231 292 261
rect 299 231 301 261
rect 42 131 44 161
rect 51 131 53 161
rect 69 131 71 161
rect 78 131 91 161
rect 98 131 118 161
rect 125 131 127 161
rect 143 131 148 161
rect 155 131 157 161
rect 173 131 175 161
rect 182 131 188 161
rect 204 131 206 161
rect 213 131 215 161
rect 260 131 262 161
rect 269 131 271 161
<< pdiffusion >>
rect 42 583 44 631
rect 51 583 53 631
rect 69 583 71 631
rect 78 583 91 631
rect 98 583 118 631
rect 125 583 127 631
rect 143 583 148 631
rect 155 583 157 631
rect 173 583 175 631
rect 182 583 188 631
rect 204 583 206 631
rect 213 583 215 631
rect 277 584 279 632
rect 286 584 288 632
rect 42 456 44 504
rect 51 456 53 504
rect 69 456 71 504
rect 78 456 91 504
rect 98 456 100 504
rect 116 456 118 504
rect 125 456 127 504
rect 204 456 206 504
rect 213 456 215 504
rect 290 456 292 504
rect 299 456 301 504
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 174 86
rect 190 76 202 86
rect 218 76 230 86
rect 246 76 258 86
rect 274 76 286 86
rect 302 76 314 86
rect 330 76 360 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
rect 50 736 62 746
rect 78 736 90 746
rect 106 736 118 746
rect 134 736 146 746
rect 162 736 174 746
rect 190 736 202 746
rect 218 736 230 746
rect 246 736 258 746
rect 274 736 286 746
rect 302 736 314 746
rect 330 736 360 746
<< ntransistor >>
rect 44 231 51 261
rect 71 231 78 261
rect 91 231 98 261
rect 118 231 125 261
rect 206 231 213 261
rect 292 231 299 261
rect 44 131 51 161
rect 71 131 78 161
rect 91 131 98 161
rect 118 131 125 161
rect 148 131 155 161
rect 175 131 182 161
rect 206 131 213 161
rect 262 131 269 161
<< ptransistor >>
rect 44 583 51 631
rect 71 583 78 631
rect 91 583 98 631
rect 118 583 125 631
rect 148 583 155 631
rect 175 583 182 631
rect 206 583 213 631
rect 279 584 286 632
rect 44 456 51 504
rect 71 456 78 504
rect 91 456 98 504
rect 118 456 125 504
rect 206 456 213 504
rect 292 456 299 504
<< polycontact >>
rect 87 695 103 711
rect 202 695 218 711
rect 49 672 73 688
rect 113 672 129 688
rect 166 672 182 688
rect 143 271 159 287
rect 253 537 269 553
rect 288 271 304 287
rect 253 191 269 207
<< ndiffcontact >>
rect 26 231 42 261
rect 53 231 69 261
rect 100 231 116 261
rect 127 231 143 261
rect 188 231 204 261
rect 215 231 231 261
rect 274 231 290 261
rect 301 231 317 261
rect 26 131 42 161
rect 53 131 69 161
rect 127 131 143 161
rect 157 131 173 161
rect 188 131 204 161
rect 215 131 231 161
rect 244 131 260 161
rect 271 131 287 161
<< pdiffcontact >>
rect 26 583 42 631
rect 53 583 69 631
rect 127 583 143 631
rect 157 583 173 631
rect 188 583 204 631
rect 215 583 231 631
rect 261 584 277 632
rect 288 584 304 632
rect 26 456 42 504
rect 53 456 69 504
rect 100 456 116 504
rect 127 456 143 504
rect 188 456 204 504
rect 215 456 231 504
rect 274 456 290 504
rect 301 456 317 504
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
rect 174 76 190 92
rect 202 76 218 92
rect 230 76 246 92
rect 258 76 274 92
rect 286 76 302 92
rect 314 76 330 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
rect 62 730 78 746
rect 90 730 106 746
rect 118 730 134 746
rect 146 730 162 746
rect 174 730 190 746
rect 202 730 218 746
rect 230 730 246 746
rect 258 730 274 746
rect 286 730 302 746
rect 314 730 330 746
<< metal1 >>
rect 0 782 360 792
rect 0 759 360 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 62 746
rect 78 730 90 746
rect 106 730 118 746
rect 134 730 146 746
rect 162 730 174 746
rect 190 730 202 746
rect 218 730 230 746
rect 246 730 258 746
rect 274 730 286 746
rect 302 730 314 746
rect 330 730 360 746
rect 0 721 360 730
rect 29 631 39 721
rect 49 688 63 697
rect 103 698 139 708
rect 153 698 202 708
rect 129 675 142 685
rect 156 675 166 685
rect 56 641 228 651
rect 56 631 66 641
rect 160 631 170 641
rect 218 631 228 641
rect 29 504 39 583
rect 129 553 141 583
rect 191 573 201 583
rect 241 573 251 721
rect 264 632 274 669
rect 294 632 304 721
rect 191 563 251 573
rect 129 541 253 553
rect 291 524 301 584
rect 56 514 140 524
rect 56 504 66 514
rect 130 504 140 514
rect 280 514 301 524
rect 280 504 290 514
rect 143 475 188 485
rect 231 474 274 484
rect 103 281 113 456
rect 317 288 327 466
rect 6 271 66 281
rect 6 101 16 271
rect 56 261 66 271
rect 103 271 143 281
rect 159 271 288 281
rect 103 261 113 271
rect 143 242 188 252
rect 231 241 274 251
rect 317 251 327 274
rect 29 221 39 231
rect 130 221 140 231
rect 29 211 140 221
rect 56 191 253 201
rect 56 161 66 191
rect 107 171 170 181
rect 29 121 39 131
rect 107 121 117 171
rect 160 161 170 171
rect 191 161 201 191
rect 279 181 289 231
rect 277 171 289 181
rect 244 161 257 167
rect 277 161 287 171
rect 29 111 117 121
rect 130 101 140 131
rect 160 121 170 131
rect 218 121 228 131
rect 160 111 228 121
rect 274 101 284 131
rect 0 92 360 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 174 92
rect 190 76 202 92
rect 218 76 230 92
rect 246 76 258 92
rect 274 76 286 92
rect 302 76 314 92
rect 330 76 360 92
rect 0 53 360 63
rect 0 30 360 40
rect 0 7 360 17
<< m2contact >>
rect 49 697 63 711
rect 139 697 153 711
rect 142 673 156 687
rect 262 669 276 683
rect 316 274 330 288
rect 241 167 255 181
<< metal2 >>
rect 48 711 60 799
rect 120 711 132 799
rect 48 697 49 711
rect 120 697 139 711
rect 48 0 60 697
rect 120 0 132 697
rect 168 687 180 799
rect 156 673 180 687
rect 168 0 180 673
rect 240 682 252 799
rect 240 670 262 682
rect 240 181 252 670
rect 312 288 324 799
rect 312 274 316 288
rect 240 167 241 181
rect 240 0 252 167
rect 312 0 324 274
<< labels >>
rlabel metal1 360 53 360 63 7 Clock
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 360 76 360 101 7 GND!
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 360 30 360 40 7 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal2 48 0 60 0 1 A
rlabel metal2 120 0 132 0 1 B
rlabel metal2 168 0 180 0 1 Cin
rlabel metal2 312 0 324 0 1 Cout
rlabel metal2 240 0 252 0 1 S
rlabel metal1 360 7 360 17 8 nReset
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 360 759 360 769 7 Scan
rlabel metal2 168 799 180 799 5 Cin
rlabel metal2 120 799 132 799 5 B
rlabel metal2 48 799 60 799 5 A
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal2 240 799 252 799 5 S
rlabel metal2 312 799 324 799 5 Cout
rlabel metal1 360 782 360 792 7 ScanReturn
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 360 721 360 746 7 Vdd!
<< end >>
