magic
tech c035u
timestamp 1386086759
<< nwell >>
rect 0 401 624 799
<< pwell >>
rect 0 0 624 401
<< polysilicon >>
rect 29 691 36 699
rect 59 691 66 699
rect 88 691 95 699
rect 115 691 122 699
rect 146 691 153 699
rect 255 691 262 719
rect 285 691 292 719
rect 336 704 403 711
rect 29 612 36 643
rect 59 599 66 643
rect 29 347 36 564
rect 59 347 66 583
rect 88 573 95 643
rect 115 591 122 643
rect 146 633 153 643
rect 149 617 153 633
rect 115 575 116 591
rect 88 347 95 557
rect 115 347 122 575
rect 146 393 153 617
rect 222 610 229 621
rect 148 377 153 393
rect 222 388 229 562
rect 255 486 262 643
rect 285 612 292 643
rect 338 612 345 623
rect 379 612 386 645
rect 396 624 403 704
rect 441 691 448 719
rect 499 691 506 719
rect 441 624 448 643
rect 396 617 448 624
rect 441 612 448 617
rect 285 486 292 564
rect 338 486 345 564
rect 379 486 386 564
rect 441 486 448 564
rect 499 532 506 643
rect 567 612 574 675
rect 29 282 36 317
rect 59 278 66 317
rect 88 309 95 317
rect 115 309 122 317
rect 146 282 153 377
rect 29 242 36 252
rect 146 244 153 252
rect 29 226 37 242
rect 222 220 229 372
rect 255 331 262 438
rect 285 402 292 438
rect 338 428 345 438
rect 354 412 366 419
rect 285 395 326 402
rect 319 358 326 395
rect 359 358 366 412
rect 379 410 386 438
rect 441 428 448 438
rect 379 403 407 410
rect 400 358 407 403
rect 441 358 448 412
rect 255 288 262 315
rect 319 288 326 328
rect 222 182 229 190
rect 255 161 262 258
rect 319 220 326 258
rect 359 220 366 328
rect 400 220 407 328
rect 441 255 448 328
rect 441 248 455 255
rect 441 225 455 232
rect 441 220 448 225
rect 499 220 506 516
rect 531 486 538 539
rect 531 358 538 438
rect 531 288 538 328
rect 255 110 262 131
rect 319 127 326 190
rect 359 128 366 190
rect 400 161 407 190
rect 441 161 448 190
rect 499 180 506 190
rect 499 142 506 150
rect 531 142 538 258
rect 567 227 574 564
rect 557 220 574 227
rect 564 190 571 195
rect 557 188 571 190
rect 564 180 571 188
rect 564 142 571 150
rect 400 120 407 131
rect 441 120 448 131
<< ndiffusion >>
rect 27 317 29 347
rect 36 317 38 347
rect 54 317 59 347
rect 66 317 88 347
rect 95 317 97 347
rect 113 317 115 347
rect 122 317 124 347
rect 27 252 29 282
rect 36 252 38 282
rect 144 252 146 282
rect 153 252 155 282
rect 314 328 319 358
rect 326 328 359 358
rect 366 328 373 358
rect 389 328 400 358
rect 407 328 441 358
rect 448 328 453 358
rect 250 258 255 288
rect 262 258 319 288
rect 326 258 337 288
rect 220 190 222 220
rect 229 190 234 220
rect 529 258 531 288
rect 538 258 544 288
rect 317 190 319 220
rect 326 190 359 220
rect 366 190 369 220
rect 433 190 441 220
rect 448 190 499 220
rect 506 190 510 220
rect 250 131 255 161
rect 262 131 267 161
rect 398 131 400 161
rect 407 131 441 161
rect 448 131 452 161
rect 561 150 564 180
rect 571 150 574 180
<< pdiffusion >>
rect 27 643 29 691
rect 36 643 38 691
rect 54 643 59 691
rect 66 643 68 691
rect 84 643 88 691
rect 95 643 97 691
rect 113 643 115 691
rect 122 643 125 691
rect 141 643 146 691
rect 153 643 156 691
rect 253 643 255 691
rect 262 643 264 691
rect 280 643 285 691
rect 292 643 294 691
rect 27 564 29 612
rect 36 564 38 612
rect 219 562 222 610
rect 229 562 234 610
rect 424 643 441 691
rect 448 643 458 691
rect 474 643 499 691
rect 506 643 509 691
rect 283 564 285 612
rect 292 564 320 612
rect 336 564 338 612
rect 345 564 355 612
rect 371 564 379 612
rect 386 564 388 612
rect 404 564 441 612
rect 448 564 450 612
rect 564 564 567 612
rect 574 564 584 612
rect 253 438 255 486
rect 262 438 265 486
rect 281 438 285 486
rect 292 438 294 486
rect 314 438 338 486
rect 345 438 353 486
rect 371 438 379 486
rect 386 438 388 486
rect 404 438 441 486
rect 448 438 451 486
rect 528 438 531 486
rect 538 438 544 486
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 198 86
rect 0 76 198 79
rect 214 76 226 86
rect 242 76 254 86
rect 270 76 282 86
rect 298 76 310 86
rect 326 76 338 86
rect 354 76 366 86
rect 382 76 394 86
rect 410 76 422 86
rect 439 76 451 86
rect 467 76 479 86
rect 495 76 507 86
rect 523 76 535 86
rect 552 76 564 86
rect 581 76 593 86
rect 610 76 624 86
<< nohmic >>
rect 0 743 198 746
rect 0 736 8 743
rect 24 736 36 743
rect 52 736 64 743
rect 80 736 92 743
rect 108 736 120 743
rect 136 736 148 743
rect 164 736 198 743
rect 214 736 226 746
rect 242 736 254 746
rect 270 736 282 746
rect 298 736 310 746
rect 326 736 338 746
rect 354 736 366 746
rect 382 736 394 746
rect 410 736 422 746
rect 438 736 450 746
rect 466 736 478 746
rect 494 736 506 746
rect 522 736 534 746
rect 550 736 562 746
rect 578 736 590 746
rect 606 736 624 746
<< ntransistor >>
rect 29 317 36 347
rect 59 317 66 347
rect 88 317 95 347
rect 115 317 122 347
rect 29 252 36 282
rect 146 252 153 282
rect 319 328 326 358
rect 359 328 366 358
rect 400 328 407 358
rect 441 328 448 358
rect 255 258 262 288
rect 319 258 326 288
rect 222 190 229 220
rect 531 258 538 288
rect 319 190 326 220
rect 359 190 366 220
rect 441 190 448 220
rect 499 190 506 220
rect 255 131 262 161
rect 400 131 407 161
rect 441 131 448 161
rect 564 150 571 180
<< ptransistor >>
rect 29 643 36 691
rect 59 643 66 691
rect 88 643 95 691
rect 115 643 122 691
rect 146 643 153 691
rect 255 643 262 691
rect 285 643 292 691
rect 29 564 36 612
rect 222 562 229 610
rect 441 643 448 691
rect 499 643 506 691
rect 285 564 292 612
rect 338 564 345 612
rect 379 564 386 612
rect 441 564 448 612
rect 567 564 574 612
rect 255 438 262 486
rect 285 438 292 486
rect 338 438 345 486
rect 379 438 386 486
rect 441 438 448 486
rect 531 438 538 486
<< polycontact >>
rect 320 695 336 711
rect 370 645 386 661
rect 59 583 75 599
rect 133 617 149 633
rect 116 575 132 591
rect 84 557 100 573
rect 132 377 148 393
rect 558 675 574 691
rect 522 539 538 555
rect 494 516 510 532
rect 213 372 229 388
rect 59 262 75 278
rect 37 226 53 242
rect 338 412 354 428
rect 441 412 457 428
rect 251 315 267 331
rect 443 232 459 248
rect 522 328 538 358
rect 391 190 407 220
rect 499 150 515 180
rect 548 190 564 220
rect 314 111 330 127
rect 355 111 372 128
<< ndiffcontact >>
rect 11 317 27 347
rect 38 317 54 347
rect 97 317 113 347
rect 124 317 140 347
rect 11 252 27 282
rect 38 252 54 282
rect 128 252 144 282
rect 155 252 175 282
rect 298 328 314 358
rect 373 328 389 358
rect 453 328 469 358
rect 234 258 250 288
rect 337 258 353 288
rect 204 190 220 220
rect 234 190 250 220
rect 513 258 529 288
rect 544 258 560 288
rect 301 190 317 220
rect 369 190 385 220
rect 417 190 433 220
rect 510 190 526 220
rect 234 131 250 161
rect 267 131 283 161
rect 382 131 398 161
rect 452 131 468 161
rect 545 150 561 180
rect 574 150 590 180
<< pdiffcontact >>
rect 11 643 27 691
rect 38 643 54 691
rect 68 643 84 691
rect 97 643 113 691
rect 125 643 141 691
rect 156 643 176 691
rect 237 643 253 691
rect 264 643 280 691
rect 294 643 310 691
rect 11 564 27 612
rect 38 564 54 612
rect 203 562 219 610
rect 234 562 250 610
rect 408 643 424 691
rect 458 643 474 691
rect 509 643 525 691
rect 267 564 283 612
rect 320 564 336 612
rect 355 564 371 612
rect 388 564 404 612
rect 450 564 466 612
rect 548 564 564 612
rect 584 564 600 612
rect 237 438 253 486
rect 265 438 281 486
rect 294 438 314 486
rect 353 438 371 486
rect 388 438 404 486
rect 451 438 467 486
rect 512 438 528 486
rect 544 438 561 486
<< psubstratetap >>
rect 6 79 22 95
rect 34 79 50 95
rect 62 79 78 95
rect 90 79 106 95
rect 118 79 134 95
rect 146 79 162 95
rect 198 76 214 92
rect 226 76 242 92
rect 254 76 270 92
rect 282 76 298 92
rect 310 76 326 92
rect 338 76 354 92
rect 366 76 382 92
rect 394 76 410 92
rect 422 76 439 92
rect 451 76 467 92
rect 479 76 495 92
rect 507 76 523 92
rect 535 76 552 92
rect 564 76 581 92
rect 593 76 610 92
<< nsubstratetap >>
rect 8 727 24 743
rect 36 727 52 743
rect 64 727 80 743
rect 92 727 108 743
rect 120 727 136 743
rect 148 727 164 743
rect 198 730 214 746
rect 226 730 242 746
rect 254 730 270 746
rect 282 730 298 746
rect 310 730 326 746
rect 338 730 354 746
rect 366 730 382 746
rect 394 730 410 746
rect 422 730 438 746
rect 450 730 466 746
rect 478 730 494 746
rect 506 730 522 746
rect 534 730 550 746
rect 562 730 578 746
rect 590 730 606 746
<< metal1 >>
rect 0 782 624 792
rect 0 759 118 769
rect 192 759 502 769
rect 518 759 624 769
rect 0 743 198 746
rect 0 727 8 743
rect 24 727 36 743
rect 52 727 64 743
rect 80 727 92 743
rect 108 727 120 743
rect 136 727 148 743
rect 164 730 198 743
rect 214 730 226 746
rect 242 730 254 746
rect 270 730 282 746
rect 298 730 310 746
rect 326 730 338 746
rect 354 730 366 746
rect 382 730 394 746
rect 410 730 422 746
rect 438 730 450 746
rect 466 730 478 746
rect 494 730 506 746
rect 522 730 534 746
rect 550 730 562 746
rect 578 730 590 746
rect 606 730 624 746
rect 164 727 624 730
rect 0 721 624 727
rect 11 691 27 721
rect 41 701 110 711
rect 41 691 51 701
rect 100 691 110 701
rect 125 691 141 721
rect 11 612 27 643
rect 71 629 81 643
rect 71 619 133 629
rect 54 583 59 599
rect 41 380 132 390
rect 41 347 51 380
rect 159 385 169 643
rect 203 634 219 721
rect 237 691 253 721
rect 264 701 320 711
rect 264 691 280 701
rect 458 701 558 711
rect 458 691 474 701
rect 558 691 574 695
rect 203 633 220 634
rect 294 633 310 643
rect 203 621 310 633
rect 320 645 370 655
rect 203 610 219 621
rect 267 612 283 621
rect 203 511 219 562
rect 320 612 336 645
rect 408 633 424 643
rect 509 633 525 643
rect 584 633 600 721
rect 355 623 600 633
rect 355 612 371 623
rect 450 612 466 623
rect 584 612 600 623
rect 234 549 250 562
rect 320 549 336 564
rect 234 539 336 549
rect 388 554 404 564
rect 388 544 522 554
rect 294 516 454 526
rect 470 516 494 526
rect 548 526 564 564
rect 510 516 564 526
rect 203 501 281 511
rect 265 486 281 501
rect 294 486 314 516
rect 584 506 600 564
rect 353 496 467 506
rect 353 486 371 496
rect 451 486 467 496
rect 512 496 600 506
rect 512 486 528 496
rect 467 438 512 486
rect 237 428 253 438
rect 388 428 404 438
rect 544 428 561 438
rect 237 418 338 428
rect 354 418 404 428
rect 457 418 561 428
rect 252 390 389 402
rect 159 375 213 385
rect 73 357 137 367
rect 14 307 24 317
rect 73 307 83 357
rect 127 347 137 357
rect 14 297 83 307
rect 54 262 59 278
rect 11 101 27 252
rect 97 101 113 317
rect 159 282 169 375
rect 252 353 265 390
rect 373 358 389 390
rect 204 341 265 353
rect 204 288 220 341
rect 251 314 267 315
rect 469 328 522 358
rect 298 318 314 328
rect 298 308 590 318
rect 204 258 234 288
rect 353 278 513 288
rect 128 101 144 252
rect 204 220 220 258
rect 234 247 250 258
rect 544 248 560 258
rect 234 235 433 247
rect 417 220 433 235
rect 459 232 560 248
rect 250 190 301 220
rect 385 190 391 220
rect 526 190 548 220
rect 204 161 220 190
rect 574 180 590 308
rect 204 131 234 161
rect 283 151 382 161
rect 515 150 545 180
rect 204 101 222 131
rect 313 111 314 127
rect 452 121 468 131
rect 372 111 468 121
rect 0 95 624 101
rect 0 79 6 95
rect 22 79 34 95
rect 50 79 62 95
rect 78 79 90 95
rect 106 79 118 95
rect 134 79 146 95
rect 162 92 624 95
rect 162 79 198 92
rect 0 76 198 79
rect 214 76 226 92
rect 242 76 254 92
rect 270 76 282 92
rect 298 76 310 92
rect 326 76 338 92
rect 354 76 366 92
rect 382 76 394 92
rect 410 76 422 92
rect 439 76 451 92
rect 467 76 479 92
rect 495 76 507 92
rect 523 76 535 92
rect 552 76 564 92
rect 581 76 593 92
rect 610 76 624 92
rect 0 53 251 63
rect 267 53 624 63
rect 0 30 39 40
rect 53 30 624 40
rect 0 7 297 17
rect 313 7 624 17
<< m2contact >>
rect 118 757 132 771
rect 502 756 518 772
rect 118 591 132 605
rect 85 543 99 557
rect 558 695 574 711
rect 454 516 470 532
rect 39 212 53 226
rect 251 298 267 314
rect 297 111 313 127
rect 251 50 267 66
rect 39 28 53 42
rect 297 3 313 19
<< metal2 >>
rect 96 557 108 799
rect 119 605 131 757
rect 99 543 108 557
rect 40 42 52 212
rect 96 0 108 543
rect 456 532 468 799
rect 504 772 516 799
rect 504 711 516 756
rect 504 695 558 711
rect 251 66 267 298
rect 297 19 313 111
rect 456 0 468 516
rect 504 0 516 695
<< labels >>
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal2 96 799 108 799 5 D
rlabel metal1 0 76 0 101 1 GND!
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 3 Clock
rlabel metal2 96 0 108 0 1 D
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal2 456 799 468 799 5 nQ
rlabel metal2 456 0 468 0 1 nQ
rlabel metal2 504 799 516 799 5 Q
rlabel metal2 504 0 516 0 1 Q
rlabel metal1 624 782 624 792 7 ScanReturn
rlabel metal1 624 759 624 769 7 Q
rlabel metal1 624 76 624 101 7 GND!
rlabel metal1 624 53 624 63 7 Clock
rlabel metal1 624 30 624 40 7 Test
rlabel metal1 624 7 624 17 7 nReset
<< end >>
