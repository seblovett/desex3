magic
tech c035u
timestamp 1385033720
<< error_ps >>
rect 1546 131 1547 132
<< metal1 >>
rect 236 906 2681 916
rect 2695 906 2797 916
rect 2811 906 2913 916
rect 1499 852 1614 862
rect 3006 852 3096 862
rect 1499 829 1614 839
rect 3006 829 3096 839
rect 1499 791 1614 816
rect 3006 791 3096 816
rect 1499 156 1614 181
rect 3006 156 3096 181
rect 1499 133 1546 143
rect 1560 133 1614 143
rect 3006 133 3096 143
rect 1499 110 1523 120
rect 1537 110 1614 120
rect 3006 110 3096 120
rect 1513 87 1614 97
rect 3006 87 3096 97
rect 1560 48 1637 58
rect 1651 48 1753 58
rect 1767 48 1870 58
rect 1537 26 1985 36
rect 1999 26 2101 36
rect 2115 26 2217 36
rect 1514 2 2333 12
rect 2347 2 2449 12
rect 2463 2 2565 12
<< m2contact >>
rect 222 905 236 919
rect 2681 904 2695 918
rect 2797 904 2811 918
rect 2913 904 2927 918
rect 1546 131 1560 145
rect 1523 108 1537 122
rect 1499 85 1513 99
rect 1546 48 1560 62
rect 1637 46 1651 60
rect 1753 46 1767 60
rect 1870 46 1884 60
rect 1523 24 1537 38
rect 1985 24 1999 38
rect 2101 24 2115 38
rect 2217 24 2231 38
rect 1500 0 1514 14
rect 2333 0 2347 14
rect 2449 0 2463 14
rect 2565 0 2579 14
<< metal2 >>
rect 223 919 235 932
rect 223 870 235 905
rect 2682 867 2694 904
rect 2798 867 2810 904
rect 2914 867 2926 904
rect 0 0 200 80
rect 223 0 235 80
rect 247 0 259 80
rect 271 0 283 80
rect 295 0 307 80
rect 1501 14 1513 85
rect 1524 38 1536 108
rect 1547 62 1559 131
rect 1638 60 1650 82
rect 1754 60 1766 82
rect 1870 60 1882 82
rect 1986 38 1998 82
rect 2102 38 2114 82
rect 2218 38 2230 82
rect 2334 14 2346 82
rect 2450 14 2462 82
rect 2566 14 2578 82
use leftbuf leftbuf_0
timestamp 1385033586
transform 1 0 -28 0 1 72
box 28 8 1527 798
use inv inv_0
timestamp 1385031732
transform 1 0 1614 0 1 82
box 0 0 116 785
use inv inv_1
timestamp 1385031732
transform 1 0 1730 0 1 82
box 0 0 116 785
use inv inv_2
timestamp 1385031732
transform 1 0 1846 0 1 82
box 0 0 116 785
use inv inv_3
timestamp 1385031732
transform 1 0 1962 0 1 82
box 0 0 116 785
use inv inv_4
timestamp 1385031732
transform 1 0 2078 0 1 82
box 0 0 116 785
use inv inv_5
timestamp 1385031732
transform 1 0 2194 0 1 82
box 0 0 116 785
use inv inv_6
timestamp 1385031732
transform 1 0 2310 0 1 82
box 0 0 116 785
use inv inv_7
timestamp 1385031732
transform 1 0 2426 0 1 82
box 0 0 116 785
use inv inv_8
timestamp 1385031732
transform 1 0 2542 0 1 82
box 0 0 116 785
use inv inv_9
timestamp 1385031732
transform 1 0 2658 0 1 82
box 0 0 116 785
use inv inv_10
timestamp 1385031732
transform 1 0 2774 0 1 82
box 0 0 116 785
use inv inv_11
timestamp 1385031732
transform 1 0 2890 0 1 82
box 0 0 116 785
<< labels >>
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 247 0 259 0 1 Test
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 295 0 307 0 1 nReset
rlabel metal2 223 932 235 932 5 SDO
rlabel metal1 3096 852 3096 862 7 nSDO
rlabel metal1 3096 829 3096 839 7 SDI
rlabel metal1 3096 791 3096 816 7 Vdd!
rlabel metal1 3096 87 3096 97 7 nResetOut
rlabel metal1 3096 110 3096 120 7 TestOut
rlabel metal1 3096 133 3096 143 7 ClockOut
rlabel metal1 3096 156 3096 181 7 GND!
<< end >>
