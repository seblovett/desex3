magic
tech c035u
timestamp 1385928100
<< metal1 >>
rect 88 803 122 813
rect 136 803 241 813
<< m2contact >>
rect 74 803 88 817
rect 122 802 136 816
rect 241 802 255 816
<< metal2 >>
rect 27 799 39 837
rect 51 799 63 837
rect 75 817 87 837
rect 75 799 87 803
rect 123 799 135 802
rect 171 799 183 837
rect 243 799 255 802
rect 291 799 303 837
use nand2 nand2_0
timestamp 1385631319
transform 1 0 3 0 1 0
box 0 0 96 799
use ../inv/inv inv_0
timestamp 1385924870
transform 1 0 99 0 1 0
box 0 0 120 799
use ../inv/inv inv_1
timestamp 1385924870
transform 1 0 219 0 1 0
box 0 0 120 799
<< labels >>
rlabel metal2 27 837 39 837 5 A
rlabel metal2 51 837 63 837 5 B
rlabel metal2 75 837 87 837 5 out
rlabel metal2 171 837 183 837 5 n1
rlabel metal2 291 837 303 837 5 n2
<< end >>
