magic
tech c035u
timestamp 1384953685
<< nwell >>
rect 0 322 281 613
<< polysilicon >>
rect 216 502 221 518
rect 28 492 35 500
rect 58 492 65 500
rect 88 492 95 500
rect 132 492 139 500
rect 162 492 169 500
rect 189 492 196 500
rect 216 492 223 502
rect 28 290 35 444
rect 58 374 65 444
rect 88 360 95 444
rect 132 374 139 444
rect 88 344 93 360
rect 58 296 65 326
rect 28 154 35 274
rect 58 250 65 280
rect 88 250 95 344
rect 132 296 139 326
rect 162 296 169 444
rect 189 322 196 444
rect 132 250 139 280
rect 88 234 93 250
rect 58 154 65 224
rect 88 154 95 234
rect 132 154 139 224
rect 162 154 169 280
rect 189 270 196 306
rect 189 154 196 254
rect 216 154 223 444
rect 246 404 251 420
rect 246 374 253 404
rect 246 250 253 326
rect 246 194 253 224
rect 251 178 253 194
rect 28 120 35 128
rect 58 120 65 128
rect 88 120 95 128
rect 132 120 139 128
rect 162 120 169 128
rect 189 120 196 128
rect 216 120 223 128
<< ndiffusion >>
rect 56 224 58 250
rect 65 224 67 250
rect 130 224 132 250
rect 139 224 141 250
rect 244 224 246 250
rect 253 224 255 250
rect 26 128 28 154
rect 35 128 58 154
rect 65 128 67 154
rect 83 128 88 154
rect 95 128 114 154
rect 130 128 132 154
rect 139 128 162 154
rect 169 128 171 154
rect 187 128 189 154
rect 196 128 216 154
rect 223 128 225 154
<< pdiffusion >>
rect 26 444 28 492
rect 35 444 40 492
rect 56 444 58 492
rect 65 444 67 492
rect 83 444 88 492
rect 95 444 114 492
rect 130 444 132 492
rect 139 444 141 492
rect 157 444 162 492
rect 169 444 171 492
rect 187 444 189 492
rect 196 444 198 492
rect 214 444 216 492
rect 223 444 225 492
rect 56 326 58 374
rect 65 326 67 374
rect 130 326 132 374
rect 139 326 141 374
rect 244 326 246 374
rect 253 326 255 374
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 174 86
rect 190 76 202 86
rect 218 76 230 86
rect 246 76 258 86
rect 274 76 281 86
rect 0 73 281 76
<< nohmic >>
rect 0 564 281 567
rect 0 557 6 564
rect 22 557 34 564
rect 50 557 62 564
rect 78 557 90 564
rect 106 557 118 564
rect 134 557 146 564
rect 162 557 174 564
rect 190 557 202 564
rect 218 557 230 564
rect 246 557 258 564
rect 274 557 281 564
<< ntransistor >>
rect 58 224 65 250
rect 132 224 139 250
rect 246 224 253 250
rect 28 128 35 154
rect 58 128 65 154
rect 88 128 95 154
rect 132 128 139 154
rect 162 128 169 154
rect 189 128 196 154
rect 216 128 223 154
<< ptransistor >>
rect 28 444 35 492
rect 58 444 65 492
rect 88 444 95 492
rect 132 444 139 492
rect 162 444 169 492
rect 189 444 196 492
rect 216 444 223 492
rect 58 326 65 374
rect 132 326 139 374
rect 246 326 253 374
<< polycontact >>
rect 221 502 237 518
rect 93 344 109 360
rect 24 274 40 290
rect 54 280 70 296
rect 180 306 196 322
rect 127 280 143 296
rect 158 280 174 296
rect 93 234 109 250
rect 180 254 196 270
rect 251 404 267 420
rect 235 178 251 194
<< ndiffcontact >>
rect 40 224 56 250
rect 67 224 83 250
rect 114 224 130 250
rect 141 224 157 250
rect 228 224 244 250
rect 255 224 271 250
rect 10 128 26 154
rect 67 128 83 154
rect 114 128 130 154
rect 171 128 187 154
rect 225 128 241 154
<< pdiffcontact >>
rect 9 444 26 492
rect 40 444 56 492
rect 67 444 83 492
rect 114 444 130 492
rect 141 444 157 492
rect 171 444 187 492
rect 198 444 214 492
rect 225 444 241 492
rect 40 326 56 374
rect 67 326 83 374
rect 114 326 130 374
rect 141 326 157 374
rect 228 326 244 374
rect 255 326 271 374
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
rect 174 76 190 92
rect 202 76 218 92
rect 230 76 246 92
rect 258 76 274 92
<< nsubstratetap >>
rect 6 548 22 564
rect 34 548 50 564
rect 62 548 78 564
rect 90 548 106 564
rect 118 548 134 564
rect 146 548 162 564
rect 174 548 190 564
rect 202 548 218 564
rect 230 548 246 564
rect 258 548 274 564
<< metal1 >>
rect 0 603 281 613
rect 0 580 174 590
rect 252 580 281 590
rect 0 564 281 567
rect 0 548 6 564
rect 22 548 34 564
rect 50 548 62 564
rect 78 548 90 564
rect 106 548 118 564
rect 134 548 146 564
rect 162 548 174 564
rect 190 548 202 564
rect 218 548 230 564
rect 246 548 258 564
rect 274 548 281 564
rect 0 542 281 548
rect 9 492 26 542
rect 67 492 83 542
rect 93 522 211 532
rect 15 394 26 444
rect 43 434 53 444
rect 93 434 103 522
rect 120 502 184 512
rect 120 492 130 502
rect 174 492 184 502
rect 201 492 211 522
rect 43 424 103 434
rect 144 414 154 444
rect 174 434 184 444
rect 228 434 238 444
rect 174 424 238 434
rect 144 404 251 414
rect 15 384 238 394
rect 40 374 50 384
rect 145 374 157 384
rect 109 344 114 360
rect 228 374 238 384
rect 73 316 83 326
rect 73 306 180 316
rect 261 305 271 326
rect 70 282 72 296
rect 120 280 127 294
rect 261 295 281 305
rect 73 260 180 270
rect 73 250 83 260
rect 261 250 271 295
rect 109 234 114 250
rect 46 214 56 224
rect 147 214 157 224
rect 228 214 238 224
rect 46 204 271 214
rect 13 184 235 194
rect 13 154 23 184
rect 70 164 150 174
rect 70 154 80 164
rect 114 98 130 128
rect 140 118 150 164
rect 174 154 184 184
rect 228 118 238 128
rect 140 108 238 118
rect 261 98 271 204
rect 0 92 281 98
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 174 92
rect 190 76 202 92
rect 218 76 230 92
rect 246 76 258 92
rect 274 76 281 92
rect 0 73 281 76
rect 0 50 281 60
rect 0 27 106 37
rect 120 27 281 37
rect 0 4 281 14
<< m2contact >>
rect 174 578 188 592
rect 238 579 252 593
rect 237 504 251 518
rect 72 282 87 296
rect 106 280 120 294
rect 174 282 188 296
rect 24 260 38 274
rect 106 25 120 39
<< metal2 >>
rect 24 274 36 617
rect 75 296 87 617
rect 175 564 187 578
rect 174 548 187 564
rect 175 296 187 548
rect 239 518 251 579
rect 24 0 36 260
rect 75 0 87 282
rect 107 39 119 280
<< labels >>
rlabel metal1 0 73 0 98 3 GND!
rlabel metal1 0 27 0 37 3 Test
rlabel metal1 0 4 0 14 2 nReset
rlabel metal1 0 50 0 60 3 Clock
rlabel metal2 24 0 36 0 1 D
rlabel metal2 75 0 87 0 1 Load
rlabel metal1 281 50 281 60 7 Clock
rlabel metal1 281 27 281 37 7 Test
rlabel metal1 281 4 281 14 8 nReset
rlabel metal1 281 73 281 98 7 GND!
rlabel metal1 281 295 281 305 7 M
rlabel metal1 281 542 281 567 1 Vdd!
rlabel metal1 281 580 281 590 7 Q
rlabel metal1 281 603 281 613 7 ScanReturn
rlabel metal1 0 603 0 613 3 ScanReturn
rlabel metal1 0 580 0 590 3 SDI
rlabel metal2 75 617 87 617 5 Load
rlabel metal2 24 617 36 617 5 D
rlabel metal1 0 542 0 567 3 Vdd!
<< end >>
