magic
tech c035u
timestamp 1385506709
<< nwell >>
rect 0 406 264 750
<< polysilicon >>
rect 24 689 31 697
rect 51 689 58 715
rect 147 689 154 697
rect 177 689 184 697
rect 232 689 239 697
rect 24 611 31 641
rect 51 611 58 641
rect 106 611 113 657
rect 24 190 31 563
rect 51 190 58 563
rect 106 190 113 563
rect 147 553 154 641
rect 177 611 184 641
rect 232 581 239 641
rect 238 565 239 581
rect 147 216 154 537
rect 177 268 184 563
rect 24 130 31 160
rect 51 130 58 160
rect 106 150 113 160
rect 147 130 154 200
rect 177 190 184 252
rect 232 206 239 565
rect 177 130 184 160
rect 232 130 239 190
rect 24 92 31 100
rect 51 92 58 100
rect 147 92 154 100
rect 177 92 184 100
rect 232 92 239 100
<< ndiffusion >>
rect 22 160 24 190
rect 31 160 51 190
rect 58 160 60 190
rect 104 160 106 190
rect 113 160 115 190
rect 175 160 177 190
rect 184 160 186 190
rect 22 100 24 130
rect 31 100 33 130
rect 49 100 51 130
rect 58 100 60 130
rect 145 100 147 130
rect 154 100 177 130
rect 184 100 186 130
rect 230 100 232 130
rect 239 100 241 130
<< pdiffusion >>
rect 22 641 24 689
rect 31 641 51 689
rect 58 641 60 689
rect 145 641 147 689
rect 154 641 159 689
rect 175 641 177 689
rect 184 641 186 689
rect 202 641 232 689
rect 239 641 241 689
rect 22 563 24 611
rect 31 563 33 611
rect 49 563 51 611
rect 58 563 60 611
rect 76 563 106 611
rect 113 563 115 611
rect 175 563 177 611
rect 184 563 186 611
<< pohmic >>
rect 0 65 6 75
rect 22 65 34 75
rect 50 65 62 75
rect 78 65 90 75
rect 106 65 118 75
rect 134 65 146 75
rect 162 65 174 75
rect 190 65 202 75
rect 218 65 230 75
rect 246 65 264 75
<< nohmic >>
rect 0 740 6 750
rect 22 740 34 750
rect 50 740 62 750
rect 78 740 90 750
rect 106 740 118 750
rect 134 740 146 750
rect 162 740 174 750
rect 190 740 202 750
rect 218 740 230 750
rect 246 740 264 750
<< ntransistor >>
rect 24 160 31 190
rect 51 160 58 190
rect 106 160 113 190
rect 177 160 184 190
rect 24 100 31 130
rect 51 100 58 130
rect 147 100 154 130
rect 177 100 184 130
rect 232 100 239 130
<< ptransistor >>
rect 24 641 31 689
rect 51 641 58 689
rect 147 641 154 689
rect 177 641 184 689
rect 232 641 239 689
rect 24 563 31 611
rect 51 563 58 611
rect 106 563 113 611
rect 177 563 184 611
<< polycontact >>
rect 101 657 117 673
rect 222 565 238 581
rect 138 537 154 553
rect 168 252 184 268
rect 138 200 154 216
rect 101 134 117 150
rect 223 190 239 206
<< ndiffcontact >>
rect 6 160 22 190
rect 60 160 76 190
rect 88 160 104 190
rect 115 160 131 190
rect 159 160 175 190
rect 186 160 202 190
rect 6 100 22 130
rect 33 100 49 130
rect 60 100 76 130
rect 129 100 145 130
rect 186 100 202 130
rect 214 100 230 130
rect 241 100 257 130
<< pdiffcontact >>
rect 6 641 22 689
rect 60 641 76 689
rect 129 641 145 689
rect 159 641 175 689
rect 186 641 202 689
rect 241 641 257 689
rect 6 563 22 611
rect 33 563 49 611
rect 60 563 76 611
rect 115 563 131 611
rect 159 563 175 611
rect 186 563 202 611
<< psubstratetap >>
rect 6 65 22 81
rect 34 65 50 81
rect 62 65 78 81
rect 90 65 106 81
rect 118 65 134 81
rect 146 65 162 81
rect 174 65 190 81
rect 202 65 218 81
rect 230 65 246 81
<< nsubstratetap >>
rect 6 734 22 750
rect 34 734 50 750
rect 62 734 78 750
rect 90 734 106 750
rect 118 734 134 750
rect 146 734 162 750
rect 174 734 190 750
rect 202 734 218 750
rect 230 734 246 750
<< metal1 >>
rect 0 780 264 790
rect 0 760 264 770
rect 0 734 6 750
rect 22 734 34 750
rect 50 734 62 750
rect 78 734 90 750
rect 106 734 118 750
rect 134 734 146 750
rect 162 734 174 750
rect 190 734 202 750
rect 218 734 230 750
rect 246 734 264 750
rect 0 725 264 734
rect 9 689 19 725
rect 132 689 142 725
rect 189 689 199 725
rect 76 660 101 670
rect 9 631 19 641
rect 135 631 145 641
rect 162 631 172 641
rect 9 621 73 631
rect 135 621 152 631
rect 162 621 231 631
rect 9 611 19 621
rect 63 611 73 621
rect 142 611 152 621
rect 142 601 159 611
rect 221 581 231 621
rect 243 605 253 641
rect 221 565 222 581
rect 36 265 46 563
rect 118 550 128 563
rect 192 553 202 563
rect 118 539 138 550
rect 36 255 168 265
rect 63 190 73 255
rect 91 206 138 216
rect 91 190 101 206
rect 192 190 202 216
rect 131 170 159 180
rect 9 130 19 160
rect 36 140 101 150
rect 36 130 46 140
rect 131 130 141 170
rect 222 190 223 206
rect 222 150 232 190
rect 189 140 232 150
rect 189 130 199 140
rect 244 130 254 166
rect 9 90 19 100
rect 63 90 73 100
rect 132 90 142 100
rect 217 90 227 100
rect 0 81 264 90
rect 0 65 6 81
rect 22 65 34 81
rect 50 65 62 81
rect 78 65 90 81
rect 106 65 118 81
rect 134 65 146 81
rect 162 65 174 81
rect 190 65 202 81
rect 218 65 230 81
rect 246 65 264 81
rect 0 45 264 55
rect 0 25 264 35
rect 0 5 264 15
<< m2contact >>
rect 47 701 61 715
rect 241 591 255 605
rect 191 539 205 553
rect 24 206 38 220
rect 191 216 205 230
rect 242 166 256 180
<< metal2 >>
rect 24 220 36 795
rect 48 715 60 795
rect 24 0 36 206
rect 48 0 60 701
rect 192 553 204 795
rect 240 605 252 795
rect 240 591 241 605
rect 192 230 204 539
rect 192 0 204 216
rect 240 180 252 591
rect 240 166 242 180
rect 240 0 252 166
<< labels >>
rlabel metal1 0 65 0 90 3 GND!
rlabel metal1 0 45 0 55 3 Clock
rlabel metal1 0 25 0 35 3 Test
rlabel metal1 0 5 0 15 3 Reset
rlabel metal2 24 0 36 0 1 A
rlabel metal2 48 0 60 0 1 B
rlabel metal2 192 0 204 0 1 C
rlabel metal2 240 0 252 0 1 S
rlabel metal2 240 795 252 795 5 S
rlabel metal2 192 795 204 795 5 C
rlabel metal2 48 795 60 795 5 B
rlabel metal2 24 795 36 795 5 A
rlabel metal1 0 780 0 790 3 ScanReturn
rlabel metal1 0 760 0 770 3 Q
rlabel metal1 0 725 0 750 3 Vdd!
rlabel metal1 264 5 264 15 7 Reset
rlabel metal1 264 25 264 35 7 Test
rlabel metal1 264 45 264 55 7 Clock
rlabel metal1 264 65 264 90 7 GND!
rlabel metal1 264 725 264 750 7 Vdd!
rlabel metal1 264 760 264 770 7 Q
rlabel metal1 264 780 264 790 7 ScanReturn
<< end >>
