magic
tech c035u
timestamp 1386086500
<< nwell >>
rect 0 401 312 799
<< pwell >>
rect 0 0 312 401
<< polysilicon >>
rect 75 697 82 711
rect 48 669 55 677
rect 75 669 82 681
rect 171 669 178 677
rect 201 669 208 677
rect 256 669 263 677
rect 48 591 55 621
rect 75 591 82 621
rect 130 591 137 637
rect 48 287 55 543
rect 50 269 55 287
rect 48 239 55 269
rect 75 239 82 543
rect 48 141 55 209
rect 75 141 82 209
rect 130 201 137 543
rect 171 533 178 621
rect 201 591 208 621
rect 256 561 263 621
rect 262 545 263 561
rect 171 227 178 517
rect 201 279 208 543
rect 130 161 137 171
rect 171 141 178 211
rect 201 201 208 263
rect 256 217 263 545
rect 201 141 208 171
rect 256 141 263 201
rect 48 103 55 111
rect 75 103 82 111
rect 171 103 178 111
rect 201 103 208 111
rect 256 103 263 111
<< ndiffusion >>
rect 46 209 48 239
rect 55 209 75 239
rect 82 209 84 239
rect 128 171 130 201
rect 137 171 139 201
rect 199 171 201 201
rect 208 171 210 201
rect 46 111 48 141
rect 55 111 57 141
rect 73 111 75 141
rect 82 111 84 141
rect 169 111 171 141
rect 178 111 201 141
rect 208 111 210 141
rect 254 111 256 141
rect 263 111 265 141
<< pdiffusion >>
rect 46 621 48 669
rect 55 621 75 669
rect 82 621 84 669
rect 169 621 171 669
rect 178 621 183 669
rect 199 621 201 669
rect 208 621 210 669
rect 226 621 256 669
rect 263 621 265 669
rect 46 543 48 591
rect 55 543 57 591
rect 73 543 75 591
rect 82 543 84 591
rect 100 543 130 591
rect 137 543 139 591
rect 199 543 201 591
rect 208 543 210 591
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 174 86
rect 190 76 202 86
rect 218 76 230 86
rect 246 76 258 86
rect 274 76 286 86
rect 302 76 312 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
rect 50 736 62 746
rect 78 736 90 746
rect 106 736 118 746
rect 134 736 146 746
rect 162 736 174 746
rect 190 736 202 746
rect 218 736 230 746
rect 246 736 258 746
rect 274 736 286 746
rect 302 736 312 746
<< ntransistor >>
rect 48 209 55 239
rect 75 209 82 239
rect 130 171 137 201
rect 201 171 208 201
rect 48 111 55 141
rect 75 111 82 141
rect 171 111 178 141
rect 201 111 208 141
rect 256 111 263 141
<< ptransistor >>
rect 48 621 55 669
rect 75 621 82 669
rect 171 621 178 669
rect 201 621 208 669
rect 256 621 263 669
rect 48 543 55 591
rect 75 543 82 591
rect 130 543 137 591
rect 201 543 208 591
<< polycontact >>
rect 71 681 87 697
rect 125 637 141 653
rect 32 269 50 287
rect 246 545 262 561
rect 162 517 178 533
rect 192 263 208 279
rect 162 211 178 227
rect 125 145 141 161
rect 247 201 263 217
<< ndiffcontact >>
rect 30 209 46 239
rect 84 209 100 239
rect 112 171 128 201
rect 139 171 155 201
rect 183 171 199 201
rect 210 171 226 201
rect 30 111 46 141
rect 57 111 73 141
rect 84 111 100 141
rect 153 111 169 141
rect 210 111 226 141
rect 238 111 254 141
rect 265 111 281 141
<< pdiffcontact >>
rect 30 621 46 669
rect 84 621 100 669
rect 153 621 169 669
rect 183 621 199 669
rect 210 621 226 669
rect 265 621 281 669
rect 30 543 46 591
rect 57 543 73 591
rect 84 543 100 591
rect 139 543 155 591
rect 183 543 199 591
rect 210 543 226 591
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
rect 174 76 190 92
rect 202 76 218 92
rect 230 76 246 92
rect 258 76 274 92
rect 286 76 302 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
rect 62 730 78 746
rect 90 730 106 746
rect 118 730 134 746
rect 146 730 162 746
rect 174 730 190 746
rect 202 730 218 746
rect 230 730 246 746
rect 258 730 274 746
rect 286 730 302 746
<< metal1 >>
rect 0 782 312 792
rect 0 759 312 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 62 746
rect 78 730 90 746
rect 106 730 118 746
rect 134 730 146 746
rect 162 730 174 746
rect 190 730 202 746
rect 218 730 230 746
rect 246 730 258 746
rect 274 730 286 746
rect 302 730 312 746
rect 0 721 312 730
rect 33 669 43 721
rect 156 669 166 721
rect 213 669 223 721
rect 100 640 125 650
rect 33 611 43 621
rect 159 611 169 621
rect 186 611 196 621
rect 33 601 97 611
rect 159 601 176 611
rect 186 601 255 611
rect 33 591 43 601
rect 87 591 97 601
rect 166 591 176 601
rect 166 581 183 591
rect 245 561 255 601
rect 267 585 277 621
rect 245 545 246 561
rect 60 276 70 543
rect 142 530 152 543
rect 216 533 226 543
rect 142 519 162 530
rect 87 276 97 291
rect 60 266 192 276
rect 87 239 97 266
rect 115 217 162 227
rect 33 141 43 209
rect 115 201 125 217
rect 216 201 226 227
rect 155 181 183 191
rect 60 151 125 161
rect 60 141 70 151
rect 155 141 165 181
rect 246 201 247 217
rect 246 161 256 201
rect 213 151 256 161
rect 213 141 223 151
rect 268 141 278 177
rect 33 101 43 111
rect 87 101 97 111
rect 156 101 166 111
rect 241 101 251 111
rect 0 92 312 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 174 92
rect 190 76 202 92
rect 218 76 230 92
rect 246 76 258 92
rect 274 76 286 92
rect 302 76 312 92
rect 0 53 312 63
rect 0 30 312 40
rect 0 7 312 17
<< m2contact >>
rect 71 697 85 711
rect 265 571 279 585
rect 36 255 50 269
rect 215 519 229 533
rect 215 227 229 241
rect 266 177 280 191
<< metal2 >>
rect 48 269 60 799
rect 72 711 84 799
rect 50 255 60 269
rect 48 0 60 255
rect 72 0 84 697
rect 216 533 228 799
rect 264 585 276 799
rect 264 571 265 585
rect 216 241 228 519
rect 216 0 228 227
rect 264 191 276 571
rect 264 177 266 191
rect 264 0 276 177
<< labels >>
rlabel metal2 48 0 60 0 1 A
rlabel metal2 72 0 84 0 1 B
rlabel metal2 216 0 228 0 1 C
rlabel metal2 264 0 276 0 1 S
rlabel metal2 264 799 276 799 5 S
rlabel metal2 216 799 228 799 5 C
rlabel metal2 72 799 84 799 5 B
rlabel metal2 48 799 60 799 5 A
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 3 nReset
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 312 76 312 101 7 GND!
rlabel metal1 312 53 312 63 7 Clock
rlabel metal1 312 30 312 40 7 Test
rlabel metal1 312 7 312 17 7 nReset
rlabel metal1 312 721 312 746 7 Vdd!
rlabel metal1 312 759 312 769 7 Scan
rlabel metal1 312 782 312 792 7 ScanReturn
<< end >>
