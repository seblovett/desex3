magic
tech c035u
timestamp 1384893035
<< nwell >>
rect 324 213 1929 425
<< polysilicon >>
rect 433 390 440 398
rect 928 390 935 398
rect 1417 390 1424 398
rect 378 291 385 299
rect 488 374 495 382
rect 515 374 522 382
rect 542 374 549 382
rect 597 378 604 386
rect 624 378 631 386
rect 651 378 658 386
rect 678 378 685 386
rect 705 378 712 386
rect 732 378 739 386
rect 759 378 766 386
rect 786 378 793 386
rect 873 291 880 299
rect 983 374 990 382
rect 1010 374 1017 382
rect 1037 374 1044 382
rect 1092 378 1099 386
rect 1119 378 1126 386
rect 1146 378 1153 386
rect 1173 378 1180 386
rect 1200 378 1207 386
rect 1227 378 1234 386
rect 1254 378 1261 386
rect 1281 378 1288 386
rect 1362 291 1369 299
rect 1472 374 1479 382
rect 1499 374 1506 382
rect 1526 374 1533 382
rect 1581 378 1588 386
rect 1608 378 1615 386
rect 1635 378 1642 386
rect 1662 378 1669 386
rect 1689 378 1696 386
rect 1716 378 1723 386
rect 1743 378 1750 386
rect 1770 378 1777 386
rect 1869 354 1871 370
rect 1864 281 1871 354
rect 378 219 385 233
rect 433 219 440 233
rect 488 219 495 233
rect 383 203 385 219
rect 438 203 440 219
rect 493 214 495 219
rect 515 214 522 233
rect 542 214 549 233
rect 597 219 604 233
rect 493 207 549 214
rect 493 203 495 207
rect 378 193 385 203
rect 433 193 440 203
rect 488 193 495 203
rect 515 193 522 207
rect 602 214 604 219
rect 624 214 631 233
rect 651 214 658 233
rect 678 214 685 233
rect 705 214 712 233
rect 732 214 739 233
rect 759 214 766 233
rect 786 216 793 233
rect 873 219 880 233
rect 928 219 935 233
rect 983 219 990 233
rect 784 214 793 216
rect 602 207 793 214
rect 602 203 604 207
rect 597 193 604 203
rect 624 193 631 207
rect 651 193 658 207
rect 678 193 685 207
rect 705 193 712 207
rect 732 193 739 207
rect 759 193 766 207
rect 786 193 793 207
rect 878 203 880 219
rect 933 203 935 219
rect 988 214 990 219
rect 1010 214 1017 233
rect 1037 214 1044 233
rect 1092 219 1099 233
rect 988 207 1044 214
rect 988 203 990 207
rect 873 193 880 203
rect 928 193 935 203
rect 983 193 990 203
rect 1010 193 1017 207
rect 1097 214 1099 219
rect 1119 214 1126 233
rect 1146 214 1153 233
rect 1173 214 1180 233
rect 1200 214 1207 233
rect 1227 214 1234 233
rect 1254 214 1261 233
rect 1281 216 1288 233
rect 1362 219 1369 233
rect 1417 219 1424 233
rect 1472 219 1479 233
rect 1279 214 1288 216
rect 1097 207 1288 214
rect 1097 203 1099 207
rect 1092 193 1099 203
rect 1119 193 1126 207
rect 1146 193 1153 207
rect 1173 193 1180 207
rect 1200 193 1207 207
rect 1227 193 1234 207
rect 1254 193 1261 207
rect 1281 193 1288 207
rect 1367 203 1369 219
rect 1422 203 1424 219
rect 1477 214 1479 219
rect 1499 214 1506 233
rect 1526 214 1533 233
rect 1581 219 1588 233
rect 1477 207 1533 214
rect 1477 203 1479 207
rect 1362 193 1369 203
rect 1417 193 1424 203
rect 1472 193 1479 203
rect 1499 193 1506 207
rect 1586 214 1588 219
rect 1608 214 1615 233
rect 1635 214 1642 233
rect 1662 214 1669 233
rect 1689 214 1696 233
rect 1716 214 1723 233
rect 1743 214 1750 233
rect 1770 216 1777 233
rect 1768 214 1777 216
rect 1586 207 1777 214
rect 1586 203 1588 207
rect 1581 193 1588 203
rect 1608 193 1615 207
rect 1635 193 1642 207
rect 1662 193 1669 207
rect 1689 193 1696 207
rect 1716 193 1723 207
rect 1743 193 1750 207
rect 1770 193 1777 207
rect 1864 193 1871 233
rect 378 165 385 173
rect 433 131 440 139
rect 873 165 880 173
rect 597 135 604 143
rect 624 135 631 143
rect 651 135 658 143
rect 678 135 685 143
rect 705 135 712 143
rect 732 135 739 143
rect 759 135 766 143
rect 786 135 793 143
rect 928 131 935 139
rect 1362 165 1369 173
rect 1092 135 1099 143
rect 1119 135 1126 143
rect 1146 135 1153 143
rect 1173 135 1180 143
rect 1200 135 1207 143
rect 1227 135 1234 143
rect 1254 135 1261 143
rect 1281 135 1288 143
rect 1417 131 1424 139
rect 1864 155 1871 163
rect 1581 135 1588 143
rect 1608 135 1615 143
rect 1635 135 1642 143
rect 1662 135 1669 143
rect 1689 135 1696 143
rect 1716 135 1723 143
rect 1743 135 1750 143
rect 1770 135 1777 143
rect 488 112 495 120
rect 515 112 522 120
rect 983 112 990 120
rect 1010 112 1017 120
rect 1472 112 1479 120
rect 1499 112 1506 120
<< ndiffusion >>
rect 376 173 378 193
rect 385 173 387 193
rect 431 139 433 193
rect 440 139 442 193
rect 486 120 488 193
rect 495 120 497 193
rect 513 120 515 193
rect 522 120 524 193
rect 595 143 597 193
rect 604 143 606 193
rect 622 143 624 193
rect 631 143 633 193
rect 649 143 651 193
rect 658 143 660 193
rect 676 143 678 193
rect 685 143 687 193
rect 703 143 705 193
rect 712 143 714 193
rect 730 143 732 193
rect 739 143 741 193
rect 757 143 759 193
rect 766 143 768 193
rect 784 143 786 193
rect 793 143 795 193
rect 871 173 873 193
rect 880 173 882 193
rect 926 139 928 193
rect 935 139 937 193
rect 981 120 983 193
rect 990 120 992 193
rect 1008 120 1010 193
rect 1017 120 1019 193
rect 1090 143 1092 193
rect 1099 143 1101 193
rect 1117 143 1119 193
rect 1126 143 1128 193
rect 1144 143 1146 193
rect 1153 143 1155 193
rect 1171 143 1173 193
rect 1180 143 1182 193
rect 1198 143 1200 193
rect 1207 143 1209 193
rect 1225 143 1227 193
rect 1234 143 1236 193
rect 1252 143 1254 193
rect 1261 143 1263 193
rect 1279 143 1281 193
rect 1288 143 1290 193
rect 1360 173 1362 193
rect 1369 173 1371 193
rect 1415 139 1417 193
rect 1424 139 1426 193
rect 1470 120 1472 193
rect 1479 120 1481 193
rect 1497 120 1499 193
rect 1506 120 1508 193
rect 1579 143 1581 193
rect 1588 143 1590 193
rect 1606 143 1608 193
rect 1615 143 1617 193
rect 1633 143 1635 193
rect 1642 143 1644 193
rect 1660 143 1662 193
rect 1669 143 1671 193
rect 1687 143 1689 193
rect 1696 143 1698 193
rect 1714 143 1716 193
rect 1723 143 1725 193
rect 1741 143 1743 193
rect 1750 143 1752 193
rect 1768 143 1770 193
rect 1777 143 1779 193
rect 1862 163 1864 193
rect 1871 163 1873 193
<< pdiffusion >>
rect 376 233 378 291
rect 385 233 387 291
rect 431 233 433 390
rect 440 233 442 390
rect 486 233 488 374
rect 495 233 497 374
rect 513 233 515 374
rect 522 233 524 374
rect 540 233 542 374
rect 549 233 551 374
rect 595 233 597 378
rect 604 233 606 378
rect 622 233 624 378
rect 631 233 633 378
rect 649 233 651 378
rect 658 233 660 378
rect 676 233 678 378
rect 685 233 687 378
rect 703 233 705 378
rect 712 233 714 378
rect 730 233 732 378
rect 739 233 741 378
rect 757 233 759 378
rect 766 233 768 378
rect 784 233 786 378
rect 793 233 795 378
rect 871 233 873 291
rect 880 233 882 291
rect 926 233 928 390
rect 935 233 937 390
rect 981 233 983 374
rect 990 233 992 374
rect 1008 233 1010 374
rect 1017 233 1019 374
rect 1035 233 1037 374
rect 1044 233 1046 374
rect 1090 233 1092 378
rect 1099 233 1101 378
rect 1117 233 1119 378
rect 1126 233 1128 378
rect 1144 233 1146 378
rect 1153 233 1155 378
rect 1171 233 1173 378
rect 1180 233 1182 378
rect 1198 233 1200 378
rect 1207 233 1209 378
rect 1225 233 1227 378
rect 1234 233 1236 378
rect 1252 233 1254 378
rect 1261 233 1263 378
rect 1279 233 1281 378
rect 1288 233 1290 378
rect 1360 233 1362 291
rect 1369 233 1371 291
rect 1415 233 1417 390
rect 1424 233 1426 390
rect 1470 233 1472 374
rect 1479 233 1481 374
rect 1497 233 1499 374
rect 1506 233 1508 374
rect 1524 233 1526 374
rect 1533 233 1535 374
rect 1579 233 1581 378
rect 1588 233 1590 378
rect 1606 233 1608 378
rect 1615 233 1617 378
rect 1633 233 1635 378
rect 1642 233 1644 378
rect 1660 233 1662 378
rect 1669 233 1671 378
rect 1687 233 1689 378
rect 1696 233 1698 378
rect 1714 233 1716 378
rect 1723 233 1725 378
rect 1741 233 1743 378
rect 1750 233 1752 378
rect 1768 233 1770 378
rect 1777 233 1779 378
rect 1862 233 1864 281
rect 1871 233 1873 281
<< pohmic >>
rect 376 85 388 95
rect 404 85 416 95
rect 432 85 444 95
rect 460 85 472 95
rect 488 85 500 95
rect 516 85 528 95
rect 544 85 556 95
rect 572 85 584 95
rect 600 85 612 95
rect 628 85 640 95
rect 656 85 668 95
rect 684 85 696 95
rect 712 85 724 95
rect 740 85 752 95
rect 768 85 780 95
rect 796 85 808 95
rect 824 85 836 95
rect 852 85 864 95
rect 880 85 892 95
rect 908 85 920 95
rect 936 85 948 95
rect 964 85 976 95
rect 992 85 1004 95
rect 1020 85 1032 95
rect 1048 85 1060 95
rect 1076 85 1088 95
rect 1104 85 1116 95
rect 1132 85 1144 95
rect 1160 85 1172 95
rect 1188 85 1200 95
rect 1216 85 1228 95
rect 1244 85 1256 95
rect 1272 85 1284 95
rect 1300 85 1312 95
rect 1328 85 1340 95
rect 1356 85 1368 95
rect 1384 85 1396 95
rect 1412 85 1424 95
rect 1440 85 1452 95
rect 1468 85 1480 95
rect 1496 85 1508 95
rect 1524 85 1536 95
rect 1552 85 1564 95
rect 1580 85 1592 95
rect 1608 85 1620 95
rect 1636 85 1648 95
rect 1664 85 1676 95
rect 1692 85 1704 95
rect 1720 85 1732 95
rect 1748 85 1760 95
rect 1776 85 1788 95
rect 1804 85 1816 95
rect 1832 85 1844 95
rect 1860 85 1872 95
rect 1888 85 1900 95
rect 1916 85 1929 95
<< nohmic >>
rect 324 415 334 425
rect 350 415 362 425
rect 378 415 390 425
rect 406 415 418 425
rect 434 415 446 425
rect 462 415 474 425
rect 490 415 502 425
rect 518 415 530 425
rect 546 415 558 425
rect 574 415 586 425
rect 602 415 614 425
rect 630 415 642 425
rect 658 415 670 425
rect 686 415 698 425
rect 714 415 726 425
rect 742 415 754 425
rect 770 415 782 425
rect 798 415 810 425
rect 826 415 838 425
rect 854 415 866 425
rect 882 415 894 425
rect 910 415 922 425
rect 938 415 950 425
rect 966 415 978 425
rect 994 415 1006 425
rect 1022 415 1034 425
rect 1050 415 1062 425
rect 1078 415 1090 425
rect 1106 415 1118 425
rect 1134 415 1146 425
rect 1162 415 1174 425
rect 1190 415 1202 425
rect 1218 415 1230 425
rect 1246 415 1258 425
rect 1274 415 1286 425
rect 1302 415 1314 425
rect 1330 415 1342 425
rect 1358 415 1370 425
rect 1386 415 1398 425
rect 1414 415 1426 425
rect 1442 415 1454 425
rect 1470 415 1482 425
rect 1498 415 1510 425
rect 1526 415 1538 425
rect 1554 415 1566 425
rect 1582 415 1594 425
rect 1610 415 1622 425
rect 1638 415 1650 425
rect 1666 415 1678 425
rect 1694 415 1706 425
rect 1722 415 1734 425
rect 1750 415 1762 425
rect 1778 415 1790 425
rect 1806 415 1818 425
rect 1834 415 1846 425
rect 1862 415 1874 425
rect 1890 415 1902 425
rect 1918 415 1929 425
<< ntransistor >>
rect 378 173 385 193
rect 433 139 440 193
rect 488 120 495 193
rect 515 120 522 193
rect 597 143 604 193
rect 624 143 631 193
rect 651 143 658 193
rect 678 143 685 193
rect 705 143 712 193
rect 732 143 739 193
rect 759 143 766 193
rect 786 143 793 193
rect 873 173 880 193
rect 928 139 935 193
rect 983 120 990 193
rect 1010 120 1017 193
rect 1092 143 1099 193
rect 1119 143 1126 193
rect 1146 143 1153 193
rect 1173 143 1180 193
rect 1200 143 1207 193
rect 1227 143 1234 193
rect 1254 143 1261 193
rect 1281 143 1288 193
rect 1362 173 1369 193
rect 1417 139 1424 193
rect 1472 120 1479 193
rect 1499 120 1506 193
rect 1581 143 1588 193
rect 1608 143 1615 193
rect 1635 143 1642 193
rect 1662 143 1669 193
rect 1689 143 1696 193
rect 1716 143 1723 193
rect 1743 143 1750 193
rect 1770 143 1777 193
rect 1864 163 1871 193
<< ptransistor >>
rect 378 233 385 291
rect 433 233 440 390
rect 488 233 495 374
rect 515 233 522 374
rect 542 233 549 374
rect 597 233 604 378
rect 624 233 631 378
rect 651 233 658 378
rect 678 233 685 378
rect 705 233 712 378
rect 732 233 739 378
rect 759 233 766 378
rect 786 233 793 378
rect 873 233 880 291
rect 928 233 935 390
rect 983 233 990 374
rect 1010 233 1017 374
rect 1037 233 1044 374
rect 1092 233 1099 378
rect 1119 233 1126 378
rect 1146 233 1153 378
rect 1173 233 1180 378
rect 1200 233 1207 378
rect 1227 233 1234 378
rect 1254 233 1261 378
rect 1281 233 1288 378
rect 1362 233 1369 291
rect 1417 233 1424 390
rect 1472 233 1479 374
rect 1499 233 1506 374
rect 1526 233 1533 374
rect 1581 233 1588 378
rect 1608 233 1615 378
rect 1635 233 1642 378
rect 1662 233 1669 378
rect 1689 233 1696 378
rect 1716 233 1723 378
rect 1743 233 1750 378
rect 1770 233 1777 378
rect 1864 233 1871 281
<< polycontact >>
rect 1853 354 1869 370
rect 367 203 383 219
rect 422 203 438 219
rect 477 203 493 219
rect 586 203 602 219
rect 862 203 878 219
rect 917 203 933 219
rect 972 203 988 219
rect 1081 203 1097 219
rect 1351 203 1367 219
rect 1406 203 1422 219
rect 1461 203 1477 219
rect 1570 203 1586 219
<< ndiffcontact >>
rect 360 173 376 193
rect 387 173 403 193
rect 415 139 431 193
rect 442 139 458 193
rect 470 120 486 193
rect 497 120 513 193
rect 524 120 540 193
rect 579 143 595 193
rect 606 143 622 193
rect 633 143 649 193
rect 660 143 676 193
rect 687 143 703 193
rect 714 143 730 193
rect 741 143 757 193
rect 768 143 784 193
rect 795 143 811 193
rect 855 173 871 193
rect 882 173 898 193
rect 910 139 926 193
rect 937 139 953 193
rect 965 120 981 193
rect 992 120 1008 193
rect 1019 120 1035 193
rect 1074 143 1090 193
rect 1101 143 1117 193
rect 1128 143 1144 193
rect 1155 143 1171 193
rect 1182 143 1198 193
rect 1209 143 1225 193
rect 1236 143 1252 193
rect 1263 143 1279 193
rect 1290 143 1306 193
rect 1344 173 1360 193
rect 1371 173 1387 193
rect 1399 139 1415 193
rect 1426 139 1442 193
rect 1454 120 1470 193
rect 1481 120 1497 193
rect 1508 120 1524 193
rect 1563 143 1579 193
rect 1590 143 1606 193
rect 1617 143 1633 193
rect 1644 143 1660 193
rect 1671 143 1687 193
rect 1698 143 1714 193
rect 1725 143 1741 193
rect 1752 143 1768 193
rect 1779 143 1795 193
rect 1846 163 1862 193
rect 1873 163 1889 193
<< pdiffcontact >>
rect 360 233 376 291
rect 387 233 403 291
rect 415 233 431 390
rect 442 233 458 390
rect 470 233 486 374
rect 497 233 513 374
rect 524 233 540 374
rect 551 233 567 374
rect 579 233 595 378
rect 606 233 622 378
rect 633 233 649 378
rect 660 233 676 378
rect 687 233 703 378
rect 714 233 730 378
rect 741 233 757 378
rect 768 233 784 378
rect 795 233 811 378
rect 855 233 871 291
rect 882 233 898 291
rect 910 233 926 390
rect 937 233 953 390
rect 965 233 981 374
rect 992 233 1008 374
rect 1019 233 1035 374
rect 1046 233 1062 374
rect 1074 233 1090 378
rect 1101 233 1117 378
rect 1128 233 1144 378
rect 1155 233 1171 378
rect 1182 233 1198 378
rect 1209 233 1225 378
rect 1236 233 1252 378
rect 1263 233 1279 378
rect 1290 233 1306 378
rect 1344 233 1360 291
rect 1371 233 1387 291
rect 1399 233 1415 390
rect 1426 233 1442 390
rect 1454 233 1470 374
rect 1481 233 1497 374
rect 1508 233 1524 374
rect 1535 233 1551 374
rect 1563 233 1579 378
rect 1590 233 1606 378
rect 1617 233 1633 378
rect 1644 233 1660 378
rect 1671 233 1687 378
rect 1698 233 1714 378
rect 1725 233 1741 378
rect 1752 233 1768 378
rect 1779 233 1795 378
rect 1846 233 1862 281
rect 1873 233 1889 281
<< psubstratetap >>
rect 360 85 376 101
rect 388 85 404 101
rect 416 85 432 101
rect 444 85 460 101
rect 472 85 488 101
rect 500 85 516 101
rect 528 85 544 101
rect 556 85 572 101
rect 584 85 600 101
rect 612 85 628 101
rect 640 85 656 101
rect 668 85 684 101
rect 696 85 712 101
rect 724 85 740 101
rect 752 85 768 101
rect 780 85 796 101
rect 808 85 824 101
rect 836 85 852 101
rect 864 85 880 101
rect 892 85 908 101
rect 920 85 936 101
rect 948 85 964 101
rect 976 85 992 101
rect 1004 85 1020 101
rect 1032 85 1048 101
rect 1060 85 1076 101
rect 1088 85 1104 101
rect 1116 85 1132 101
rect 1144 85 1160 101
rect 1172 85 1188 101
rect 1200 85 1216 101
rect 1228 85 1244 101
rect 1256 85 1272 101
rect 1284 85 1300 101
rect 1312 85 1328 101
rect 1340 85 1356 101
rect 1368 85 1384 101
rect 1396 85 1412 101
rect 1424 85 1440 101
rect 1452 85 1468 101
rect 1480 85 1496 101
rect 1508 85 1524 101
rect 1536 85 1552 101
rect 1564 85 1580 101
rect 1592 85 1608 101
rect 1620 85 1636 101
rect 1648 85 1664 101
rect 1676 85 1692 101
rect 1704 85 1720 101
rect 1732 85 1748 101
rect 1760 85 1776 101
rect 1788 85 1804 101
rect 1816 85 1832 101
rect 1844 85 1860 101
rect 1872 85 1888 101
rect 1900 85 1916 101
<< nsubstratetap >>
rect 334 409 350 425
rect 362 409 378 425
rect 390 409 406 425
rect 418 409 434 425
rect 446 409 462 425
rect 474 409 490 425
rect 502 409 518 425
rect 530 409 546 425
rect 558 409 574 425
rect 586 409 602 425
rect 614 409 630 425
rect 642 409 658 425
rect 670 409 686 425
rect 698 409 714 425
rect 726 409 742 425
rect 754 409 770 425
rect 782 409 798 425
rect 810 409 826 425
rect 838 409 854 425
rect 866 409 882 425
rect 894 409 910 425
rect 922 409 938 425
rect 950 409 966 425
rect 978 409 994 425
rect 1006 409 1022 425
rect 1034 409 1050 425
rect 1062 409 1078 425
rect 1090 409 1106 425
rect 1118 409 1134 425
rect 1146 409 1162 425
rect 1174 409 1190 425
rect 1202 409 1218 425
rect 1230 409 1246 425
rect 1258 409 1274 425
rect 1286 409 1302 425
rect 1314 409 1330 425
rect 1342 409 1358 425
rect 1370 409 1386 425
rect 1398 409 1414 425
rect 1426 409 1442 425
rect 1454 409 1470 425
rect 1482 409 1498 425
rect 1510 409 1526 425
rect 1538 409 1554 425
rect 1566 409 1582 425
rect 1594 409 1610 425
rect 1622 409 1638 425
rect 1650 409 1666 425
rect 1678 409 1694 425
rect 1706 409 1722 425
rect 1734 409 1750 425
rect 1762 409 1778 425
rect 1790 409 1806 425
rect 1818 409 1834 425
rect 1846 409 1862 425
rect 1874 409 1890 425
rect 1902 409 1918 425
<< metal1 >>
rect 236 463 1831 473
rect 1875 463 1929 473
rect 236 439 1929 449
rect 185 409 334 425
rect 350 409 362 425
rect 378 409 390 425
rect 406 409 418 425
rect 434 409 446 425
rect 462 409 474 425
rect 490 409 502 425
rect 518 409 530 425
rect 546 409 558 425
rect 574 409 586 425
rect 602 409 614 425
rect 630 409 642 425
rect 658 409 670 425
rect 686 409 698 425
rect 714 409 726 425
rect 742 409 754 425
rect 770 409 782 425
rect 798 409 810 425
rect 826 409 838 425
rect 854 409 866 425
rect 882 409 894 425
rect 910 409 922 425
rect 938 409 950 425
rect 966 409 978 425
rect 994 409 1006 425
rect 1022 409 1034 425
rect 1050 409 1062 425
rect 1078 409 1090 425
rect 1106 409 1118 425
rect 1134 409 1146 425
rect 1162 409 1174 425
rect 1190 409 1202 425
rect 1218 409 1230 425
rect 1246 409 1258 425
rect 1274 409 1286 425
rect 1302 409 1314 425
rect 1330 409 1342 425
rect 1358 409 1370 425
rect 1386 409 1398 425
rect 1414 409 1426 425
rect 1442 409 1454 425
rect 1470 409 1482 425
rect 1498 409 1510 425
rect 1526 409 1538 425
rect 1554 409 1566 425
rect 1582 409 1594 425
rect 1610 409 1622 425
rect 1638 409 1650 425
rect 1666 409 1678 425
rect 1694 409 1706 425
rect 1722 409 1734 425
rect 1750 409 1762 425
rect 1778 409 1790 425
rect 1806 409 1818 425
rect 1834 409 1846 425
rect 1862 409 1874 425
rect 1890 409 1902 425
rect 1918 409 1929 425
rect 185 400 1929 409
rect 360 291 376 400
rect 415 390 431 400
rect 470 374 486 400
rect 524 374 540 400
rect 579 378 595 400
rect 633 378 649 400
rect 687 378 703 400
rect 741 378 757 400
rect 795 378 811 400
rect 855 291 871 400
rect 910 390 926 400
rect 965 374 981 400
rect 1019 374 1035 400
rect 1074 378 1090 400
rect 1128 378 1144 400
rect 1182 378 1198 400
rect 1236 378 1252 400
rect 1290 378 1306 400
rect 1344 291 1360 400
rect 1399 390 1415 400
rect 1454 374 1470 400
rect 1508 374 1524 400
rect 1563 378 1579 400
rect 1617 378 1633 400
rect 1671 378 1687 400
rect 1725 378 1741 400
rect 1779 378 1795 400
rect 1855 370 1869 376
rect 1879 281 1889 400
rect 284 204 367 214
rect 393 216 403 233
rect 393 206 422 216
rect 393 193 403 206
rect 448 216 458 233
rect 448 206 477 216
rect 448 193 458 206
rect 503 216 513 233
rect 557 216 567 233
rect 503 206 586 216
rect 503 193 513 206
rect 612 216 622 233
rect 666 216 676 233
rect 720 216 730 233
rect 774 216 784 233
rect 612 206 794 216
rect 612 193 622 206
rect 666 193 676 206
rect 720 193 730 206
rect 774 193 784 206
rect 843 207 862 217
rect 888 216 898 233
rect 888 206 917 216
rect 888 193 898 206
rect 943 216 953 233
rect 943 206 972 216
rect 943 193 953 206
rect 998 216 1008 233
rect 1052 216 1062 233
rect 998 206 1081 216
rect 998 193 1008 206
rect 1107 216 1117 233
rect 1161 216 1171 233
rect 1215 216 1225 233
rect 1269 216 1279 233
rect 1107 206 1295 216
rect 1107 193 1117 206
rect 1161 193 1171 206
rect 1215 193 1225 206
rect 1269 193 1279 206
rect 1336 205 1351 215
rect 1377 216 1387 233
rect 1377 206 1406 216
rect 1377 193 1387 206
rect 1432 216 1442 233
rect 1432 206 1461 216
rect 1432 193 1442 206
rect 1487 216 1497 233
rect 1541 216 1551 233
rect 1487 206 1570 216
rect 1487 193 1497 206
rect 1596 216 1606 233
rect 1650 216 1660 233
rect 1704 216 1714 233
rect 1758 216 1768 233
rect 1596 206 1806 216
rect 1596 193 1606 206
rect 1650 193 1660 206
rect 1704 193 1714 206
rect 1758 193 1768 206
rect 1846 193 1856 233
rect 360 110 376 173
rect 415 110 431 139
rect 470 110 486 120
rect 524 110 540 120
rect 579 110 595 143
rect 633 110 649 143
rect 687 110 703 143
rect 741 110 757 143
rect 795 110 811 143
rect 855 110 871 173
rect 910 110 926 139
rect 965 110 981 120
rect 1019 110 1035 120
rect 1074 110 1090 143
rect 1128 110 1144 143
rect 1182 110 1198 143
rect 1236 110 1252 143
rect 1290 110 1306 143
rect 1344 110 1360 173
rect 1399 110 1415 139
rect 1454 110 1470 120
rect 1508 110 1524 120
rect 1563 110 1579 143
rect 1617 110 1633 143
rect 1671 110 1687 143
rect 1725 110 1741 143
rect 1779 110 1795 143
rect 1873 110 1883 163
rect 360 101 1929 110
rect 376 85 388 101
rect 404 85 416 101
rect 432 85 444 101
rect 460 85 472 101
rect 488 85 500 101
rect 516 85 528 101
rect 544 85 556 101
rect 572 85 584 101
rect 600 85 612 101
rect 628 85 640 101
rect 656 85 668 101
rect 684 85 696 101
rect 712 85 724 101
rect 740 85 752 101
rect 768 85 780 101
rect 796 85 808 101
rect 824 85 836 101
rect 852 85 864 101
rect 880 85 892 101
rect 908 85 920 101
rect 936 85 948 101
rect 964 85 976 101
rect 992 85 1004 101
rect 1020 85 1032 101
rect 1048 85 1060 101
rect 1076 85 1088 101
rect 1104 85 1116 101
rect 1132 85 1144 101
rect 1160 85 1172 101
rect 1188 85 1200 101
rect 1216 85 1228 101
rect 1244 85 1256 101
rect 1272 85 1284 101
rect 1300 85 1312 101
rect 1328 85 1340 101
rect 1356 85 1368 101
rect 1384 85 1396 101
rect 1412 85 1424 101
rect 1440 85 1452 101
rect 1468 85 1480 101
rect 1496 85 1508 101
rect 1524 85 1536 101
rect 1552 85 1564 101
rect 1580 85 1592 101
rect 1608 85 1620 101
rect 1636 85 1648 101
rect 1664 85 1676 101
rect 1692 85 1704 101
rect 1720 85 1732 101
rect 1748 85 1760 101
rect 1776 85 1788 101
rect 1804 85 1816 101
rect 1832 85 1844 101
rect 1860 85 1872 101
rect 1888 85 1900 101
rect 1916 85 1929 101
rect 808 61 1929 71
rect 260 39 828 49
rect 1309 37 1929 47
rect 308 15 1322 25
rect 1819 13 1929 23
<< m2contact >>
rect 222 461 236 475
rect 1831 460 1845 474
rect 1861 460 1875 474
rect 222 437 236 451
rect 171 400 185 425
rect 1855 376 1869 390
rect 270 202 284 216
rect 794 203 808 217
rect 829 204 843 218
rect 1295 204 1309 218
rect 1322 204 1336 218
rect 1806 204 1820 218
rect 1832 205 1846 219
rect 794 61 808 75
rect 246 37 260 51
rect 828 37 842 51
rect 1295 35 1309 49
rect 294 13 308 27
rect 1322 12 1336 26
rect 1805 11 1819 25
<< metal2 >>
rect 0 425 200 509
rect 223 475 235 509
rect 0 400 171 425
rect 185 400 200 425
rect 0 0 200 400
rect 223 0 235 437
rect 247 51 259 509
rect 271 216 283 509
rect 247 0 259 37
rect 271 0 283 202
rect 295 27 307 509
rect 1833 219 1845 460
rect 1861 390 1873 460
rect 1869 376 1873 390
rect 795 75 807 203
rect 830 51 842 204
rect 1296 49 1308 204
rect 1323 26 1335 204
rect 1467 83 1479 103
rect 1502 83 1514 103
rect 295 0 307 13
rect 1806 25 1818 204
<< labels >>
rlabel metal2 295 509 307 509 5 nReset
rlabel metal2 271 509 283 509 5 Clock
rlabel metal2 247 509 259 509 5 Test
rlabel metal2 223 509 235 509 5 SDO
rlabel metal2 0 509 200 509 5 Vdd!
rlabel metal1 1929 400 1929 425 7 Vdd!
rlabel metal1 1929 85 1929 110 7 GND!
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 295 0 307 0 1 nReset
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 247 0 259 0 1 Test
rlabel metal1 1929 439 1929 449 7 SDI
rlabel metal1 1929 463 1929 473 7 nSDO
rlabel metal1 1929 61 1929 71 7 ClockOut
rlabel metal1 1929 37 1929 47 7 TestOut
rlabel metal1 1929 13 1929 23 7 nResetOut
<< end >>
