magic
tech c035u
timestamp 1385929574
<< error_ps >>
rect 47 834 48 835
<< metal1 >>
rect -35 860 71 870
rect -155 836 47 846
rect -275 813 24 823
rect 109 813 144 823
rect 158 813 263 823
<< m2contact >>
rect -49 860 -35 874
rect 71 858 85 872
rect -169 834 -155 848
rect 47 834 61 848
rect -289 809 -275 823
rect 24 811 38 825
rect 95 809 109 823
rect 144 811 158 825
rect 263 811 277 825
<< metal2 >>
rect -336 799 -324 891
rect -288 799 -276 809
rect -216 799 -204 891
rect -168 799 -156 834
rect -96 799 -84 891
rect -48 799 -36 860
rect 24 825 36 891
rect 48 848 60 891
rect 72 872 84 891
rect 24 799 36 811
rect 48 799 60 834
rect 72 799 84 858
rect 96 823 108 891
rect 96 799 108 809
rect 144 799 156 811
rect 192 799 204 891
rect 264 799 276 811
rect 312 799 324 891
use inv inv_2
timestamp 1385924870
transform 1 0 -360 0 1 0
box 0 0 120 799
use inv inv_3
timestamp 1385924870
transform 1 0 -240 0 1 0
box 0 0 120 799
use inv inv_4
timestamp 1385924870
transform 1 0 -120 0 1 0
box 0 0 120 799
use nand3 nand3_0
timestamp 1385920731
transform 1 0 0 0 1 0
box 0 0 120 799
use inv inv_0
timestamp 1385924870
transform 1 0 120 0 1 0
box 0 0 120 799
use inv inv_1
timestamp 1385924870
transform 1 0 240 0 1 0
box 0 0 120 799
<< labels >>
rlabel metal2 312 891 324 891 5 n2
rlabel metal2 192 891 204 891 5 n1
rlabel metal2 96 891 108 891 5 Y
rlabel metal2 72 891 84 891 5 C
rlabel metal2 48 891 60 891 5 B
rlabel metal2 24 891 36 891 5 A
rlabel metal2 -336 891 -324 891 5 NA
rlabel metal2 -216 891 -204 891 5 NB
rlabel metal2 -96 891 -84 891 5 NC
<< end >>
