magic
tech c035u
timestamp 1386235766
<< nwell >>
rect 0 401 1464 799
<< pwell >>
rect 0 0 1464 401
<< polysilicon >>
rect 538 711 545 719
rect 565 711 572 719
rect 592 711 599 719
rect 619 711 626 719
rect 875 711 882 719
rect 902 711 909 719
rect 929 711 936 719
rect 956 711 963 719
rect 1212 711 1219 719
rect 1239 711 1246 719
rect 1266 711 1273 719
rect 1293 711 1300 719
rect 480 633 487 641
rect 507 633 514 641
rect 425 578 432 586
rect 370 479 377 487
rect 817 633 824 641
rect 844 633 851 641
rect 762 578 769 586
rect 707 479 714 487
rect 1154 633 1161 641
rect 1181 633 1188 641
rect 1099 578 1106 586
rect 1044 479 1051 487
rect 1394 516 1396 532
rect 1389 471 1396 516
rect 370 388 377 421
rect 425 388 432 421
rect 480 389 487 421
rect 375 372 377 388
rect 430 372 432 388
rect 485 385 487 389
rect 507 385 514 421
rect 538 389 545 421
rect 485 378 514 385
rect 485 373 487 378
rect 543 385 545 389
rect 565 385 572 421
rect 592 385 599 421
rect 619 385 626 421
rect 707 388 714 421
rect 762 388 769 421
rect 817 389 824 421
rect 543 378 626 385
rect 543 373 545 378
rect 370 362 377 372
rect 425 362 432 372
rect 480 362 487 373
rect 538 362 545 373
rect 565 362 572 378
rect 712 372 714 388
rect 767 372 769 388
rect 822 385 824 389
rect 844 385 851 421
rect 875 389 882 421
rect 822 378 851 385
rect 822 373 824 378
rect 880 385 882 389
rect 902 385 909 421
rect 929 385 936 421
rect 956 385 963 421
rect 1044 388 1051 421
rect 1099 388 1106 421
rect 1154 389 1161 421
rect 880 378 963 385
rect 880 373 882 378
rect 707 362 714 372
rect 762 362 769 372
rect 817 362 824 373
rect 875 362 882 373
rect 902 362 909 378
rect 1049 372 1051 388
rect 1104 372 1106 388
rect 1159 385 1161 389
rect 1181 385 1188 421
rect 1212 389 1219 421
rect 1159 378 1188 385
rect 1159 373 1161 378
rect 1217 385 1219 389
rect 1239 385 1246 421
rect 1266 385 1273 421
rect 1293 385 1300 421
rect 1217 378 1300 385
rect 1217 373 1219 378
rect 1044 362 1051 372
rect 1099 362 1106 372
rect 1154 362 1161 373
rect 1212 362 1219 373
rect 1239 362 1246 378
rect 1389 377 1396 423
rect 370 334 377 342
rect 425 300 432 308
rect 480 208 487 216
rect 707 334 714 342
rect 762 300 769 308
rect 817 208 824 216
rect 1044 334 1051 342
rect 1099 300 1106 308
rect 1154 208 1161 216
rect 1389 339 1396 347
rect 538 154 545 162
rect 565 154 572 162
rect 875 154 882 162
rect 902 154 909 162
rect 1212 154 1219 162
rect 1239 154 1246 162
<< ndiffusion >>
rect 368 342 370 362
rect 377 342 379 362
rect 423 308 425 362
rect 432 308 434 362
rect 478 216 480 362
rect 487 216 489 362
rect 536 162 538 362
rect 545 162 547 362
rect 563 162 565 362
rect 572 162 574 362
rect 705 342 707 362
rect 714 342 716 362
rect 760 308 762 362
rect 769 308 771 362
rect 815 216 817 362
rect 824 216 826 362
rect 873 162 875 362
rect 882 162 884 362
rect 900 162 902 362
rect 909 162 911 362
rect 1042 342 1044 362
rect 1051 342 1053 362
rect 1097 308 1099 362
rect 1106 308 1108 362
rect 1152 216 1154 362
rect 1161 216 1163 362
rect 1210 162 1212 362
rect 1219 162 1221 362
rect 1237 162 1239 362
rect 1246 162 1248 362
rect 1387 347 1389 377
rect 1396 347 1398 377
<< pdiffusion >>
rect 368 421 370 479
rect 377 421 379 479
rect 423 421 425 578
rect 432 421 434 578
rect 478 421 480 633
rect 487 421 489 633
rect 505 421 507 633
rect 514 421 516 633
rect 536 421 538 711
rect 545 421 547 711
rect 563 421 565 711
rect 572 421 574 711
rect 590 421 592 711
rect 599 421 601 711
rect 617 421 619 711
rect 626 421 628 711
rect 705 421 707 479
rect 714 421 716 479
rect 760 421 762 578
rect 769 421 771 578
rect 815 421 817 633
rect 824 421 826 633
rect 842 421 844 633
rect 851 421 853 633
rect 873 421 875 711
rect 882 421 884 711
rect 900 421 902 711
rect 909 421 911 711
rect 927 421 929 711
rect 936 421 938 711
rect 954 421 956 711
rect 963 421 965 711
rect 1042 421 1044 479
rect 1051 421 1053 479
rect 1097 421 1099 578
rect 1106 421 1108 578
rect 1152 421 1154 633
rect 1161 421 1163 633
rect 1179 421 1181 633
rect 1188 421 1190 633
rect 1210 421 1212 711
rect 1219 421 1221 711
rect 1237 421 1239 711
rect 1246 421 1248 711
rect 1264 421 1266 711
rect 1273 421 1275 711
rect 1291 421 1293 711
rect 1300 421 1302 711
rect 1387 423 1389 471
rect 1396 423 1398 471
<< pohmic >>
rect 320 76 326 86
rect 342 76 354 86
rect 370 76 382 86
rect 398 76 410 86
rect 426 76 438 86
rect 454 76 466 86
rect 482 76 494 86
rect 510 76 522 86
rect 538 76 550 86
rect 567 76 579 86
rect 595 76 607 86
rect 623 76 635 86
rect 651 76 663 86
rect 679 76 691 86
rect 707 76 719 86
rect 735 76 747 86
rect 763 76 775 86
rect 791 76 803 86
rect 819 76 831 86
rect 847 76 859 86
rect 875 76 887 86
rect 904 76 916 86
rect 932 76 944 86
rect 960 76 972 86
rect 988 76 1000 86
rect 1016 76 1028 86
rect 1044 76 1056 86
rect 1072 76 1084 86
rect 1100 76 1112 86
rect 1128 76 1140 86
rect 1156 76 1168 86
rect 1184 76 1196 86
rect 1212 76 1224 86
rect 1241 76 1253 86
rect 1269 76 1281 86
rect 1297 76 1309 86
rect 1325 76 1337 86
rect 1353 76 1365 86
rect 1381 76 1393 86
rect 1409 76 1421 86
rect 1437 76 1464 86
<< nohmic >>
rect 202 736 214 746
rect 230 736 242 746
rect 258 736 270 746
rect 286 736 298 746
rect 314 736 326 746
rect 342 736 354 746
rect 370 736 382 746
rect 398 736 410 746
rect 426 736 438 746
rect 454 736 466 746
rect 482 736 494 746
rect 510 736 522 746
rect 538 736 550 746
rect 567 736 579 746
rect 595 736 607 746
rect 623 736 635 746
rect 651 736 663 746
rect 679 736 691 746
rect 707 736 719 746
rect 735 736 747 746
rect 763 736 775 746
rect 791 736 803 746
rect 819 736 831 746
rect 847 736 859 746
rect 875 736 887 746
rect 904 736 916 746
rect 932 736 944 746
rect 960 736 972 746
rect 988 736 1000 746
rect 1016 736 1028 746
rect 1044 736 1056 746
rect 1072 736 1084 746
rect 1100 736 1112 746
rect 1128 736 1140 746
rect 1156 736 1168 746
rect 1184 736 1196 746
rect 1212 736 1224 746
rect 1241 736 1253 746
rect 1269 736 1281 746
rect 1297 736 1309 746
rect 1325 736 1337 746
rect 1353 736 1365 746
rect 1381 736 1393 746
rect 1409 736 1421 746
rect 1437 736 1464 746
<< ntransistor >>
rect 370 342 377 362
rect 425 308 432 362
rect 480 216 487 362
rect 538 162 545 362
rect 565 162 572 362
rect 707 342 714 362
rect 762 308 769 362
rect 817 216 824 362
rect 875 162 882 362
rect 902 162 909 362
rect 1044 342 1051 362
rect 1099 308 1106 362
rect 1154 216 1161 362
rect 1212 162 1219 362
rect 1239 162 1246 362
rect 1389 347 1396 377
<< ptransistor >>
rect 370 421 377 479
rect 425 421 432 578
rect 480 421 487 633
rect 507 421 514 633
rect 538 421 545 711
rect 565 421 572 711
rect 592 421 599 711
rect 619 421 626 711
rect 707 421 714 479
rect 762 421 769 578
rect 817 421 824 633
rect 844 421 851 633
rect 875 421 882 711
rect 902 421 909 711
rect 929 421 936 711
rect 956 421 963 711
rect 1044 421 1051 479
rect 1099 421 1106 578
rect 1154 421 1161 633
rect 1181 421 1188 633
rect 1212 421 1219 711
rect 1239 421 1246 711
rect 1266 421 1273 711
rect 1293 421 1300 711
rect 1389 423 1396 471
<< polycontact >>
rect 1378 516 1394 532
rect 359 372 375 388
rect 414 372 430 388
rect 469 373 485 389
rect 527 373 543 389
rect 696 372 712 388
rect 751 372 767 388
rect 806 373 822 389
rect 864 373 880 389
rect 1033 372 1049 388
rect 1088 372 1104 388
rect 1143 373 1159 389
rect 1201 373 1217 389
<< ndiffcontact >>
rect 352 342 368 362
rect 379 342 395 362
rect 407 308 423 362
rect 434 308 450 362
rect 462 216 478 362
rect 489 216 505 362
rect 520 162 536 362
rect 547 162 563 362
rect 574 162 590 362
rect 689 342 705 362
rect 716 342 732 362
rect 744 308 760 362
rect 771 308 787 362
rect 799 216 815 362
rect 826 216 842 362
rect 857 162 873 362
rect 884 162 900 362
rect 911 162 927 362
rect 1026 342 1042 362
rect 1053 342 1069 362
rect 1081 308 1097 362
rect 1108 308 1124 362
rect 1136 216 1152 362
rect 1163 216 1179 362
rect 1194 162 1210 362
rect 1221 162 1237 362
rect 1248 162 1264 362
rect 1371 347 1387 377
rect 1398 347 1414 377
<< pdiffcontact >>
rect 519 633 536 711
rect 352 421 368 479
rect 379 421 395 479
rect 407 421 423 578
rect 434 421 450 578
rect 462 421 478 633
rect 489 421 505 633
rect 516 421 536 633
rect 547 421 563 711
rect 574 421 590 711
rect 601 421 617 711
rect 628 421 644 711
rect 856 633 873 711
rect 689 421 705 479
rect 716 421 732 479
rect 744 421 760 578
rect 771 421 787 578
rect 799 421 815 633
rect 826 421 842 633
rect 853 421 873 633
rect 884 421 900 711
rect 911 421 927 711
rect 938 421 954 711
rect 965 421 981 711
rect 1193 633 1210 711
rect 1026 421 1042 479
rect 1053 421 1069 479
rect 1081 421 1097 578
rect 1108 421 1124 578
rect 1136 421 1152 633
rect 1163 421 1179 633
rect 1190 421 1210 633
rect 1221 421 1237 711
rect 1248 421 1264 711
rect 1275 421 1291 711
rect 1302 421 1318 711
rect 1371 423 1387 471
rect 1398 423 1414 471
<< psubstratetap >>
rect 352 312 368 328
rect 407 279 423 295
rect 462 187 478 203
rect 689 313 705 329
rect 744 279 760 295
rect 799 187 815 203
rect 1026 313 1042 329
rect 1081 279 1097 295
rect 1136 187 1152 203
rect 1398 318 1414 334
rect 326 76 342 92
rect 354 76 370 92
rect 382 76 398 92
rect 410 76 426 92
rect 438 76 454 92
rect 466 76 482 92
rect 494 76 510 92
rect 522 76 538 92
rect 550 76 567 92
rect 579 76 595 92
rect 607 76 623 92
rect 635 76 651 92
rect 663 76 679 92
rect 691 76 707 92
rect 719 76 735 92
rect 747 76 763 92
rect 775 76 791 92
rect 803 76 819 92
rect 831 76 847 92
rect 859 76 875 92
rect 887 76 904 92
rect 916 76 932 92
rect 944 76 960 92
rect 972 76 988 92
rect 1000 76 1016 92
rect 1028 76 1044 92
rect 1056 76 1072 92
rect 1084 76 1100 92
rect 1112 76 1128 92
rect 1140 76 1156 92
rect 1168 76 1184 92
rect 1196 76 1212 92
rect 1224 76 1241 92
rect 1253 76 1269 92
rect 1281 76 1297 92
rect 1309 76 1325 92
rect 1337 76 1353 92
rect 1365 76 1381 92
rect 1393 76 1409 92
rect 1421 76 1437 92
<< nsubstratetap >>
rect 214 730 230 746
rect 242 730 258 746
rect 270 730 286 746
rect 298 730 314 746
rect 326 730 342 746
rect 354 730 370 746
rect 382 730 398 746
rect 410 730 426 746
rect 438 730 454 746
rect 466 730 482 746
rect 494 730 510 746
rect 522 730 538 746
rect 550 730 567 746
rect 579 730 595 746
rect 607 730 623 746
rect 635 730 651 746
rect 663 730 679 746
rect 691 730 707 746
rect 719 730 735 746
rect 747 730 763 746
rect 775 730 791 746
rect 803 730 819 746
rect 831 730 847 746
rect 859 730 875 746
rect 887 730 904 746
rect 916 730 932 746
rect 944 730 960 746
rect 972 730 988 746
rect 1000 730 1016 746
rect 1028 730 1044 746
rect 1056 730 1072 746
rect 1084 730 1100 746
rect 1112 730 1128 746
rect 1140 730 1156 746
rect 1168 730 1184 746
rect 1196 730 1212 746
rect 1224 730 1241 746
rect 1253 730 1269 746
rect 1281 730 1297 746
rect 1309 730 1325 746
rect 1337 730 1353 746
rect 1365 730 1381 746
rect 1393 730 1409 746
rect 1421 730 1437 746
<< metal1 >>
rect 185 756 200 792
rect 229 782 1356 792
rect 1395 782 1464 792
rect 229 759 1464 769
rect 200 730 214 746
rect 230 730 242 746
rect 258 730 270 746
rect 286 730 298 746
rect 314 730 326 746
rect 342 730 354 746
rect 370 730 382 746
rect 398 730 410 746
rect 426 730 438 746
rect 454 730 466 746
rect 482 730 494 746
rect 510 730 522 746
rect 538 730 550 746
rect 567 730 579 746
rect 595 730 607 746
rect 623 730 635 746
rect 651 730 663 746
rect 679 730 691 746
rect 707 730 719 746
rect 735 730 747 746
rect 763 730 775 746
rect 791 730 803 746
rect 819 730 831 746
rect 847 730 859 746
rect 875 730 887 746
rect 904 730 916 746
rect 932 730 944 746
rect 960 730 972 746
rect 988 730 1000 746
rect 1016 730 1028 746
rect 1044 730 1056 746
rect 1072 730 1084 746
rect 1100 730 1112 746
rect 1128 730 1140 746
rect 1156 730 1168 746
rect 1184 730 1196 746
rect 1212 730 1224 746
rect 1241 730 1253 746
rect 1269 730 1281 746
rect 1297 730 1309 746
rect 1325 730 1337 746
rect 1353 730 1365 746
rect 1381 730 1393 746
rect 1409 730 1421 746
rect 1437 730 1464 746
rect 200 721 1464 730
rect 352 479 368 721
rect 407 578 423 721
rect 462 633 478 721
rect 516 711 536 721
rect 574 711 590 721
rect 628 711 644 721
rect 516 633 519 711
rect 689 479 705 721
rect 744 578 760 721
rect 799 633 815 721
rect 853 711 873 721
rect 911 711 927 721
rect 965 711 981 721
rect 853 633 856 711
rect 1026 479 1042 721
rect 1081 578 1097 721
rect 1136 633 1152 721
rect 1190 711 1210 721
rect 1248 711 1264 721
rect 1302 711 1318 721
rect 1190 633 1193 711
rect 1404 471 1414 721
rect 240 349 252 387
rect 277 375 359 385
rect 263 363 277 373
rect 385 385 395 421
rect 385 375 414 385
rect 385 362 395 375
rect 440 386 450 421
rect 440 376 469 386
rect 440 362 450 376
rect 495 386 505 421
rect 495 376 527 386
rect 495 362 505 376
rect 553 387 563 421
rect 607 389 617 421
rect 553 377 606 387
rect 553 362 563 377
rect 722 385 732 421
rect 722 375 751 385
rect 722 362 732 375
rect 777 386 787 421
rect 777 376 806 386
rect 777 362 787 376
rect 832 386 842 421
rect 832 376 864 386
rect 832 362 842 376
rect 890 387 900 421
rect 944 389 954 421
rect 890 377 944 387
rect 890 362 900 377
rect 1059 385 1069 421
rect 1059 375 1088 385
rect 1059 362 1069 375
rect 1114 386 1124 421
rect 1114 376 1143 386
rect 1114 362 1124 376
rect 1169 386 1179 421
rect 1169 376 1201 386
rect 1169 362 1179 376
rect 1227 387 1237 421
rect 1281 389 1291 421
rect 1227 377 1279 387
rect 1227 362 1237 377
rect 1371 377 1381 423
rect 352 328 368 342
rect 352 101 368 312
rect 407 295 423 308
rect 407 101 423 279
rect 462 203 478 216
rect 462 101 478 187
rect 520 101 536 162
rect 574 101 590 162
rect 689 329 705 342
rect 689 101 705 313
rect 744 295 760 308
rect 744 101 760 279
rect 799 203 815 216
rect 799 101 815 187
rect 857 101 873 162
rect 911 101 927 162
rect 1026 329 1042 342
rect 1026 101 1042 313
rect 1081 295 1097 308
rect 1081 101 1097 279
rect 1136 203 1152 216
rect 1136 101 1152 187
rect 1194 101 1210 162
rect 1248 101 1264 162
rect 1398 334 1408 347
rect 1398 101 1408 318
rect 320 92 1464 101
rect 320 76 326 92
rect 342 76 354 92
rect 370 76 382 92
rect 398 76 410 92
rect 426 76 438 92
rect 454 76 466 92
rect 482 76 494 92
rect 510 76 522 92
rect 538 76 550 92
rect 567 76 579 92
rect 595 76 607 92
rect 623 76 635 92
rect 651 76 663 92
rect 679 76 691 92
rect 707 76 719 92
rect 735 76 747 92
rect 763 76 775 92
rect 791 76 803 92
rect 819 76 831 92
rect 847 76 859 92
rect 875 76 887 92
rect 904 76 916 92
rect 932 76 944 92
rect 960 76 972 92
rect 988 76 1000 92
rect 1016 76 1028 92
rect 1044 76 1056 92
rect 1072 76 1084 92
rect 1100 76 1112 92
rect 1128 76 1140 92
rect 1156 76 1168 92
rect 1184 76 1196 92
rect 1212 76 1224 92
rect 1241 76 1253 92
rect 1269 76 1281 92
rect 1297 76 1309 92
rect 1325 76 1337 92
rect 1353 76 1365 92
rect 1381 76 1393 92
rect 1409 76 1421 92
rect 1437 76 1464 92
rect 216 5 228 67
rect 239 43 253 53
rect 620 53 1464 63
rect 253 30 681 40
rect 959 30 1464 40
rect 301 7 1018 17
rect 1042 7 1270 17
rect 1294 7 1304 17
rect 1318 7 1464 17
<< m2contact >>
rect 215 780 229 794
rect 1356 781 1370 795
rect 1381 781 1395 795
rect 215 756 229 770
rect 0 721 200 746
rect 1380 532 1394 546
rect 1357 457 1371 471
rect 263 373 277 387
rect 263 349 277 363
rect 606 375 620 389
rect 682 373 696 387
rect 944 375 958 389
rect 1019 373 1033 387
rect 1279 375 1293 389
rect 239 53 253 67
rect 606 51 620 65
rect 239 29 253 43
rect 681 28 695 42
rect 945 29 959 43
rect 239 5 253 19
rect 263 5 277 19
rect 287 5 301 19
rect 1018 5 1032 19
rect 1280 5 1294 19
rect 1304 5 1318 19
<< metal2 >>
rect 0 746 200 799
rect 216 794 228 799
rect 0 0 200 721
rect 216 0 228 756
rect 240 67 252 799
rect 264 387 276 799
rect 264 363 276 373
rect 240 43 252 53
rect 240 19 252 29
rect 264 19 276 349
rect 288 19 300 799
rect 1358 471 1370 781
rect 1382 546 1394 781
rect 607 65 619 375
rect 682 42 694 373
rect 946 43 958 375
rect 1019 19 1031 373
rect 1281 19 1293 375
rect 1294 5 1304 19
rect 240 0 252 5
rect 264 0 276 5
rect 288 0 300 5
<< labels >>
rlabel metal2 0 799 200 799 5 Vdd!
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal1 1464 721 1464 746 7 Vdd!
rlabel metal1 1464 759 1464 769 7 SDI
rlabel metal1 1464 782 1464 792 7 nSDO
rlabel metal1 1464 53 1464 63 7 ClockOut
rlabel metal1 1464 30 1464 40 7 TestOut
rlabel metal1 1464 7 1464 17 7 nResetOut
rlabel metal1 1464 76 1464 101 7 GND!
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 288 799 300 799 5 nReset
rlabel metal2 240 799 252 799 5 Test
rlabel metal2 264 799 276 799 5 Clock
rlabel metal2 216 799 228 799 5 SDO
<< end >>
