* HSPICE file created from rdtype.ext - technology: c035u

.option scale=0.05u

m1000 active_100_481 Clk Vdd Vdd pmos03553 w=48 l=7
m1001 Vdd nRst active_100_481 Vdd pmos03553 w=48 l=7
m1002 active_67_416 D Vdd Vdd pmos03553 w=48 l=7
m1003 Q active_100_481 Vdd Vdd pmos03553 w=48 l=7
m1004 Vdd nQ Q Vdd pmos03553 w=48 l=7
m1005 active_67_416 nRst Vdd Vdd pmos03553 w=48 l=7
m1006 Vdd active_75_348 active_67_416 Vdd pmos03553 w=48 l=7
m1007 active_224_416 active_67_416 Vdd Vdd pmos03553 w=48 l=7
m1008 Vdd active_100_481 active_224_416 Vdd pmos03553 w=48 l=7
m1009 Vdd Clk active_75_348 Vdd pmos03553 w=48 l=7
m1010 nQ nRst Vdd Vdd pmos03553 w=48 l=7
m1011 Vdd active_75_348 nQ Vdd pmos03553 w=48 l=7
m1012 active_75_348 active_67_416 Vdd Vdd pmos03553 w=48 l=7
m1013 Vdd active_100_481 active_75_348 Vdd pmos03553 w=48 l=7
m1014 active_164_267 nRst active_136_259 GND nmos03553 w=30 l=7
m1015 GND active_75_348 active_164_267 GND nmos03553 w=30 l=7
m1016 active_245_267 active_67_416 GND GND nmos03553 w=30 l=7
m1017 active_224_416 active_100_481 active_245_267 GND nmos03553 w=30 l=7
m1018 active_100_217 Clk GND GND nmos03553 w=30 l=7
m1019 active_164_217 nRst active_100_217 GND nmos03553 w=30 l=7
m1020 active_67_169 D GND GND nmos03553 w=30 l=7
m1021 Vdd Q nQ Vdd pmos03553 w=48 l=7
m1022 active_100_481 active_224_416 Vdd Vdd pmos03553 w=48 l=7
m1023 active_100_481 active_224_416 active_164_217 GND nmos03553 w=30 l=7
m1024 active_164_169 nRst active_67_169 GND nmos03553 w=30 l=7
m1025 active_67_416 active_75_348 active_164_169 GND nmos03553 w=30 l=7
m1026 active_286_169 active_100_481 GND GND nmos03553 w=30 l=7
m1027 Q nQ active_286_169 GND nmos03553 w=30 l=7
m1028 active_100_127 Clk GND GND nmos03553 w=30 l=7
m1029 active_245_127 active_67_416 active_100_127 GND nmos03553 w=30 l=7
m1030 active_75_348 active_100_481 active_245_127 GND nmos03553 w=30 l=7
m1031 active_136_259 Q nQ GND nmos03553 w=30 l=7
C0 Test GND 2.0fF **FLOATING
C1 ScanReturn GND 2.0fF **FLOATING
C2 active_164_217 GND 0.7fF
C3 active_136_259 GND 1.8fF
C4 active_224_416 GND 2.1fF
C5 Q GND 6.7fF
C6 active_75_348 GND 2.3fF
C7 active_67_416 GND 1.9fF
C8 D GND 1.5fF
C9 nQ GND 5.6fF
C10 active_100_481 GND 3.2fF
C11 nRst GND 3.6fF
C12 Clk GND 4.3fF
C13 Vdd GND 6.1fF

** hspice subcircuit dictionary
