magic
tech c035u
timestamp 1384969111
<< nwell >>
rect 0 219 117 308
<< polysilicon >>
rect 28 274 35 282
rect 55 274 62 282
rect 82 274 89 282
rect 28 202 35 226
rect 33 186 35 202
rect 28 68 35 186
rect 55 156 62 226
rect 82 179 89 226
rect 88 163 89 179
rect 61 140 62 156
rect 55 68 62 140
rect 82 68 89 163
rect 28 30 35 38
rect 55 30 62 38
rect 82 30 89 38
<< ndiffusion >>
rect 26 38 28 68
rect 35 38 55 68
rect 62 38 64 68
rect 80 38 82 68
rect 89 38 91 68
<< pdiffusion >>
rect 26 226 28 274
rect 35 226 37 274
rect 53 226 55 274
rect 62 226 64 274
rect 80 226 82 274
rect 89 226 91 274
<< pohmic >>
rect 0 7 6 14
rect 22 7 34 14
rect 50 7 62 14
rect 78 7 90 14
rect 106 7 117 14
rect 0 4 117 7
<< nohmic >>
rect 0 305 117 308
rect 0 298 6 305
rect 22 298 34 305
rect 50 298 62 305
rect 78 298 90 305
rect 106 298 117 305
<< ntransistor >>
rect 28 38 35 68
rect 55 38 62 68
rect 82 38 89 68
<< ptransistor >>
rect 28 226 35 274
rect 55 226 62 274
rect 82 226 89 274
<< polycontact >>
rect 17 186 33 202
rect 72 163 88 179
rect 45 140 61 156
<< ndiffcontact >>
rect 10 38 26 68
rect 64 38 80 68
rect 91 38 107 68
<< pdiffcontact >>
rect 10 226 26 274
rect 37 226 53 274
rect 64 226 80 274
rect 91 226 107 274
<< psubstratetap >>
rect 6 7 22 23
rect 34 7 50 23
rect 62 7 78 23
rect 90 7 106 23
<< nsubstratetap >>
rect 6 289 22 305
rect 34 289 50 305
rect 62 289 78 305
rect 90 289 106 305
<< metal1 >>
rect 0 305 117 308
rect 0 289 6 305
rect 22 289 34 305
rect 50 289 62 305
rect 78 289 90 305
rect 106 289 117 305
rect 0 284 117 289
rect 10 274 26 284
rect 64 274 80 284
rect 107 226 108 236
rect 43 176 53 226
rect 10 166 72 176
rect 10 68 20 166
rect 98 153 108 226
rect 97 68 107 139
rect 64 28 80 38
rect 0 23 117 28
rect 0 7 6 23
rect 22 7 34 23
rect 50 7 62 23
rect 78 7 90 23
rect 106 7 117 23
rect 0 4 117 7
<< m2contact >>
rect 17 202 31 216
rect 46 126 60 140
rect 96 139 110 153
<< metal2 >>
rect 24 274 36 312
rect 24 226 37 274
rect 24 216 36 226
rect 31 202 36 216
rect 24 23 36 202
rect 48 156 60 312
rect 48 140 61 156
rect 96 153 108 312
rect 23 7 36 23
rect 24 0 36 7
rect 48 0 60 126
rect 96 0 108 139
<< labels >>
rlabel metal1 0 284 0 308 3 Vdd!
rlabel metal2 24 312 36 312 5 A
rlabel metal2 48 312 60 312 5 B
rlabel metal2 48 0 60 0 1 B
rlabel metal2 24 0 36 0 1 A
rlabel metal1 0 4 0 28 3 GND!
rlabel metal2 96 0 108 0 1 Y
rlabel metal2 96 312 108 312 5 Y
rlabel metal1 117 4 117 28 7 GND!
rlabel metal1 117 284 117 308 7 Vdd!
<< end >>
