magic
tech c035u
timestamp 1385077924
<< nwell >>
rect 0 523 100 735
<< polysilicon >>
rect 32 571 39 579
rect 59 571 66 579
rect 32 504 39 523
rect 38 488 39 504
rect 59 499 66 523
rect 32 453 39 488
rect 65 483 66 499
rect 59 453 66 483
rect 32 415 39 423
rect 59 415 66 423
<< ndiffusion >>
rect 30 423 32 453
rect 39 423 41 453
rect 57 423 59 453
rect 66 423 68 453
<< pdiffusion >>
rect 30 523 32 571
rect 39 523 59 571
rect 66 523 68 571
<< pohmic >>
rect 0 75 6 85
rect 22 75 34 85
rect 50 75 62 85
rect 78 75 100 85
<< nohmic >>
rect 0 725 6 735
rect 22 725 34 735
rect 50 725 62 735
rect 78 725 100 735
<< ntransistor >>
rect 32 423 39 453
rect 59 423 66 453
<< ptransistor >>
rect 32 523 39 571
rect 59 523 66 571
<< polycontact >>
rect 22 488 38 504
rect 49 483 65 499
<< ndiffcontact >>
rect 6 423 30 453
rect 41 423 57 453
rect 68 423 92 453
<< pdiffcontact >>
rect 6 523 30 571
rect 68 523 94 571
<< psubstratetap >>
rect 6 75 22 91
rect 34 75 50 91
rect 62 75 78 91
<< nsubstratetap >>
rect 6 719 22 735
rect 34 719 50 735
rect 62 719 78 735
<< metal1 >>
rect 0 771 100 781
rect 0 748 100 758
rect 0 719 6 735
rect 22 719 34 735
rect 50 719 62 735
rect 78 719 100 735
rect 0 710 100 719
rect 5 575 30 710
rect 6 571 30 575
rect 77 499 87 523
rect 77 473 87 485
rect 47 463 87 473
rect 47 453 57 463
rect 6 100 30 423
rect 68 100 92 423
rect 0 91 100 100
rect 0 75 6 91
rect 22 75 34 91
rect 50 75 62 91
rect 78 75 100 91
rect 0 52 100 62
rect 0 29 100 39
rect 0 6 100 16
<< m2contact >>
rect 48 499 62 513
rect 23 474 37 488
rect 75 485 89 499
<< metal2 >>
rect 24 504 36 787
rect 22 488 36 504
rect 48 513 60 787
rect 72 499 84 787
rect 24 0 36 474
rect 48 0 60 499
rect 72 485 75 499
rect 72 0 84 485
<< labels >>
rlabel metal2 24 787 36 787 5 A
rlabel metal2 24 0 36 0 1 A
rlabel metal2 48 0 60 0 1 B
rlabel metal2 48 787 60 787 5 B
rlabel metal2 72 787 84 787 5 Y
rlabel metal2 72 0 84 0 1 Y
rlabel metal1 0 710 0 735 3 Vdd!
rlabel metal1 100 710 100 735 1 Vdd!
rlabel metal1 100 748 100 758 1 Scan
rlabel metal1 100 771 100 781 1 ScanReturn
rlabel metal1 0 771 0 781 3 ScanReturn
rlabel metal1 0 748 0 758 3 Scan
rlabel metal1 0 6 0 16 3 nReset
rlabel metal1 100 6 100 16 7 nReset
rlabel metal1 100 29 100 39 7 Test
rlabel metal1 0 29 0 39 3 Test
rlabel metal1 0 52 0 62 3 Clock
rlabel metal1 100 52 100 62 7 Clock
rlabel metal1 0 75 0 100 3 GND!
rlabel metal1 100 75 100 100 7 GND!
<< end >>
