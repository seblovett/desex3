magic
tech c035u
timestamp 1385058581
<< error_s >>
rect 352 570 357 572
rect 1336 168 1337 174
<< metal1 >>
rect 236 908 2624 918
rect 2638 908 2740 918
rect 2754 908 2856 918
rect 1442 854 1557 864
rect 2949 854 3039 864
rect 1442 831 1557 841
rect 2949 831 3039 841
rect 1442 793 1557 818
rect 2949 793 3039 818
rect 1442 158 1557 183
rect 2949 158 3039 183
rect 1442 135 1509 145
rect 1523 135 1557 145
rect 2949 135 3039 145
rect 1442 112 1486 122
rect 1500 112 1557 122
rect 2949 112 3039 122
rect 1442 89 1462 99
rect 1476 89 1557 99
rect 2949 89 3039 99
rect 1523 50 1580 60
rect 1594 50 1696 60
rect 1710 50 1813 60
rect 1500 28 1928 38
rect 1942 28 2044 38
rect 2058 28 2160 38
rect 1477 4 2276 14
rect 2290 4 2392 14
rect 2406 4 2508 14
<< m2contact >>
rect 222 907 236 921
rect 2624 906 2638 920
rect 2740 906 2754 920
rect 2856 906 2870 920
rect 1509 134 1523 148
rect 1486 110 1500 124
rect 1462 87 1476 101
rect 1509 50 1523 64
rect 1580 48 1594 62
rect 1696 48 1710 62
rect 1813 48 1827 62
rect 1486 26 1500 40
rect 1928 26 1942 40
rect 2044 26 2058 40
rect 2160 26 2174 40
rect 1463 2 1477 16
rect 2276 2 2290 16
rect 2392 2 2406 16
rect 2508 2 2522 16
<< metal2 >>
rect 223 921 235 934
rect 223 872 235 907
rect 2625 869 2637 906
rect 2741 869 2753 906
rect 2857 869 2869 906
rect 0 0 200 80
rect 223 0 235 80
rect 247 0 259 80
rect 271 0 283 80
rect 295 0 307 80
rect 1464 16 1476 87
rect 1487 40 1499 110
rect 1510 64 1522 134
rect 1581 62 1593 84
rect 1697 62 1709 84
rect 1813 62 1825 84
rect 1929 40 1941 84
rect 2045 40 2057 84
rect 2161 40 2173 84
rect 2277 16 2289 84
rect 2393 16 2405 84
rect 2509 16 2521 84
use leftbuf leftbuf_0
timestamp 1385058125
transform 1 0 0 0 1 82
box 0 -2 1442 790
use inv inv_0
timestamp 1385031732
transform 1 0 1557 0 1 84
box 0 0 116 785
use inv inv_1
timestamp 1385031732
transform 1 0 1673 0 1 84
box 0 0 116 785
use inv inv_2
timestamp 1385031732
transform 1 0 1789 0 1 84
box 0 0 116 785
use inv inv_3
timestamp 1385031732
transform 1 0 1905 0 1 84
box 0 0 116 785
use inv inv_4
timestamp 1385031732
transform 1 0 2021 0 1 84
box 0 0 116 785
use inv inv_5
timestamp 1385031732
transform 1 0 2137 0 1 84
box 0 0 116 785
use inv inv_6
timestamp 1385031732
transform 1 0 2253 0 1 84
box 0 0 116 785
use inv inv_7
timestamp 1385031732
transform 1 0 2369 0 1 84
box 0 0 116 785
use inv inv_8
timestamp 1385031732
transform 1 0 2485 0 1 84
box 0 0 116 785
use inv inv_9
timestamp 1385031732
transform 1 0 2601 0 1 84
box 0 0 116 785
use inv inv_10
timestamp 1385031732
transform 1 0 2717 0 1 84
box 0 0 116 785
use inv inv_11
timestamp 1385031732
transform 1 0 2833 0 1 84
box 0 0 116 785
<< labels >>
rlabel metal1 3039 854 3039 864 7 nSDO
rlabel metal1 3039 831 3039 841 7 SDI
rlabel metal1 3039 793 3039 818 7 Vdd!
rlabel metal1 3039 89 3039 99 7 nResetOut
rlabel metal1 3039 112 3039 122 7 TestOut
rlabel metal1 3039 135 3039 145 7 ClockOut
rlabel metal1 3039 158 3039 183 7 GND!
rlabel metal2 223 934 235 934 5 SDO
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 247 0 259 0 1 Test
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 295 0 307 0 1 nReset
<< end >>
