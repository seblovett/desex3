magic
tech c035u
timestamp 1386444371
<< metal1 >>
rect 23 878 114 888
rect 23 824 33 878
rect 368 874 738 884
rect 22 814 43 824
rect 0 776 43 801
rect 835 430 876 440
rect 890 430 906 440
rect 0 131 43 156
rect 12 85 43 95
rect 12 30 22 85
rect 12 20 234 30
rect 440 24 546 35
rect 560 24 877 34
<< m2contact >>
rect 114 874 128 888
rect 354 872 368 886
rect 738 872 752 886
rect 876 428 890 442
rect 234 20 248 34
rect 426 23 440 37
rect 546 22 560 36
rect 877 24 891 38
<< metal2 >>
rect 67 854 79 913
rect 115 888 127 913
rect 115 854 127 874
rect 307 854 319 913
rect 355 854 367 872
rect 475 854 487 913
rect 595 854 607 913
rect 739 886 751 913
rect 739 854 751 872
rect 187 0 199 55
rect 235 34 247 55
rect 427 37 439 55
rect 547 36 559 55
rect 878 38 890 428
rect 235 0 247 20
use inv inv_0
timestamp 1386238110
transform 1 0 43 0 1 55
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 163 0 1 55
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 283 0 1 55
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 403 0 1 55
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 523 0 1 55
box 0 0 120 799
use smux2 smux2_0
timestamp 1386234984
transform 1 0 643 0 1 55
box 0 0 192 799
<< labels >>
rlabel metal1 0 131 0 156 3 GND!
rlabel metal1 0 776 0 801 3 Vdd!
rlabel metal1 906 430 906 440 7 M
rlabel metal2 595 913 607 913 5 n2
rlabel metal2 475 913 487 913 5 n1
rlabel metal2 739 913 751 913 5 D
rlabel metal2 307 913 319 913 5 ND
rlabel metal2 235 0 247 0 1 TEST
rlabel metal2 187 0 199 0 1 NTEST
rlabel metal2 115 913 127 913 5 SDI
rlabel metal2 67 913 79 913 5 NSDI
<< end >>
