magic
tech c035u
timestamp 1384775938
<< nwell >>
rect 0 320 281 565
<< polysilicon >>
rect 216 503 221 519
rect 28 490 35 498
rect 58 490 65 498
rect 88 490 95 498
rect 132 490 139 498
rect 162 490 169 498
rect 189 490 196 498
rect 216 490 223 503
rect 28 314 35 442
rect 58 372 65 442
rect 88 358 95 442
rect 132 372 139 442
rect 88 342 93 358
rect 28 132 35 298
rect 58 294 65 324
rect 58 228 65 278
rect 88 223 95 342
rect 132 228 139 324
rect 162 274 169 442
rect 189 320 196 442
rect 88 207 93 223
rect 58 132 65 202
rect 88 132 95 207
rect 132 132 139 202
rect 162 132 169 258
rect 189 248 196 304
rect 189 132 196 232
rect 216 132 223 442
rect 246 402 251 418
rect 246 372 253 402
rect 246 228 253 324
rect 246 172 253 202
rect 251 156 253 172
rect 28 98 35 106
rect 58 98 65 106
rect 88 98 95 106
rect 132 41 139 106
rect 162 98 169 106
rect 189 98 196 106
rect 216 98 223 106
<< ndiffusion >>
rect 56 202 58 228
rect 65 202 67 228
rect 130 202 132 228
rect 139 202 141 228
rect 244 202 246 228
rect 253 202 255 228
rect 26 106 28 132
rect 35 106 58 132
rect 65 106 67 132
rect 83 106 88 132
rect 95 106 114 132
rect 130 106 132 132
rect 139 106 162 132
rect 169 106 171 132
rect 187 106 189 132
rect 196 106 216 132
rect 223 106 225 132
<< pdiffusion >>
rect 26 442 28 490
rect 35 442 40 490
rect 56 442 58 490
rect 65 442 67 490
rect 83 442 88 490
rect 95 442 114 490
rect 130 442 132 490
rect 139 442 141 490
rect 157 442 162 490
rect 169 442 171 490
rect 187 442 189 490
rect 196 442 198 490
rect 214 442 216 490
rect 223 442 225 490
rect 56 324 58 372
rect 65 324 67 372
rect 130 324 132 372
rect 139 324 141 372
rect 244 324 246 372
rect 253 324 255 372
<< ntransistor >>
rect 58 202 65 228
rect 132 202 139 228
rect 246 202 253 228
rect 28 106 35 132
rect 58 106 65 132
rect 88 106 95 132
rect 132 106 139 132
rect 162 106 169 132
rect 189 106 196 132
rect 216 106 223 132
<< ptransistor >>
rect 28 442 35 490
rect 58 442 65 490
rect 88 442 95 490
rect 132 442 139 490
rect 162 442 169 490
rect 189 442 196 490
rect 216 442 223 490
rect 58 324 65 372
rect 132 324 139 372
rect 246 324 253 372
<< polycontact >>
rect 221 503 237 519
rect 93 342 109 358
rect 24 298 40 314
rect 54 278 70 294
rect 180 304 196 320
rect 158 258 174 274
rect 93 207 109 223
rect 180 232 196 248
rect 251 402 267 418
rect 235 156 251 172
rect 124 25 140 41
<< ndiffcontact >>
rect 40 202 56 228
rect 67 202 83 228
rect 114 202 130 228
rect 141 202 157 228
rect 228 202 244 228
rect 255 202 271 228
rect 10 106 26 132
rect 67 106 83 132
rect 114 106 130 132
rect 171 106 187 132
rect 225 106 241 132
<< pdiffcontact >>
rect 9 442 26 490
rect 40 442 56 490
rect 67 442 83 490
rect 114 442 130 490
rect 141 442 157 490
rect 171 442 187 490
rect 198 442 214 490
rect 225 442 241 490
rect 40 324 56 372
rect 67 324 83 372
rect 114 324 130 372
rect 141 324 157 372
rect 228 324 244 372
rect 255 324 271 372
<< psubstratetap >>
rect 7 54 23 70
rect 228 56 244 72
<< nsubstratetap >>
rect 7 543 23 559
rect 228 544 244 560
<< metal1 >>
rect 0 560 281 565
rect 0 559 228 560
rect 0 543 7 559
rect 23 544 228 559
rect 244 544 281 560
rect 23 543 281 544
rect 0 540 281 543
rect 9 490 26 540
rect 67 490 83 540
rect 93 520 211 530
rect 15 392 26 442
rect 43 432 53 442
rect 93 432 103 520
rect 120 500 184 510
rect 120 490 130 500
rect 174 490 184 500
rect 201 490 211 520
rect 237 505 281 515
rect 43 422 103 432
rect 144 412 154 442
rect 174 432 184 442
rect 228 432 238 442
rect 174 422 238 432
rect 144 402 251 412
rect 15 382 238 392
rect 40 372 50 382
rect 145 372 157 382
rect 109 342 114 358
rect 228 372 238 382
rect 73 314 83 324
rect 73 304 180 314
rect 24 295 38 298
rect 70 278 72 292
rect 261 283 271 324
rect 0 258 158 268
rect 261 273 281 283
rect 73 238 180 248
rect 73 228 83 238
rect 261 228 271 273
rect 109 207 114 223
rect 46 192 56 202
rect 147 192 157 202
rect 228 192 238 202
rect 46 182 271 192
rect 13 162 235 172
rect 13 132 23 162
rect 70 142 150 152
rect 70 132 80 142
rect 114 76 130 106
rect 140 96 150 142
rect 174 132 184 162
rect 228 96 238 106
rect 140 86 238 96
rect 261 76 271 182
rect 0 72 281 76
rect 0 70 228 72
rect 0 54 7 70
rect 23 56 228 70
rect 244 56 281 72
rect 23 54 281 56
rect 0 51 281 54
rect 0 31 124 41
<< m2contact >>
rect 24 281 38 295
rect 72 278 87 292
<< metal2 >>
rect 24 295 36 569
rect 75 292 87 569
rect 24 25 36 281
rect 75 25 87 278
<< labels >>
rlabel metal2 24 569 36 569 5 D
rlabel metal2 75 569 87 569 5 Load
rlabel metal1 0 540 0 565 3 Vdd!
rlabel metal1 281 505 281 515 7 Q
rlabel metal1 281 540 281 565 1 Vdd!
rlabel metal1 281 273 281 283 7 M
rlabel metal1 281 51 281 76 7 GND!
rlabel metal1 0 51 0 76 3 GND!
rlabel metal2 75 25 87 25 1 Load
rlabel metal2 24 25 36 25 1 D
rlabel metal1 0 31 0 41 3 Test
rlabel metal1 0 258 0 268 3 SDI
<< end >>
