magic
tech c035u
timestamp 1384878722
<< nwell >>
rect 32 505 439 566
rect 32 345 438 505
<< polysilicon >>
rect 93 529 100 537
rect 123 529 130 537
rect 279 529 286 537
rect 337 529 344 541
rect 169 522 241 529
rect 60 464 67 475
rect 60 304 67 416
rect 93 396 100 481
rect 123 464 130 481
rect 176 464 183 475
rect 217 464 224 480
rect 234 476 241 522
rect 279 476 286 481
rect 234 469 286 476
rect 279 464 286 469
rect 337 417 344 481
rect 405 464 412 513
rect 123 396 130 416
rect 176 396 183 416
rect 217 396 224 416
rect 279 396 286 416
rect 93 304 100 348
rect 123 319 130 348
rect 176 338 183 348
rect 192 322 204 329
rect 123 312 164 319
rect 157 297 164 312
rect 197 297 204 322
rect 217 326 224 348
rect 279 338 286 348
rect 217 319 245 326
rect 238 297 245 319
rect 279 297 286 322
rect 60 199 67 288
rect 93 247 100 288
rect 157 247 164 267
rect 60 161 67 169
rect 93 157 100 217
rect 157 199 164 217
rect 197 199 204 267
rect 238 199 245 267
rect 279 226 286 267
rect 279 210 281 226
rect 279 199 286 210
rect 337 199 344 401
rect 369 396 376 421
rect 369 297 376 348
rect 369 247 376 281
rect 157 136 164 169
rect 197 137 204 169
rect 238 157 245 169
rect 279 157 286 169
rect 337 158 344 169
rect 93 119 100 127
rect 238 119 245 127
rect 279 119 286 127
rect 337 120 344 128
rect 369 120 376 217
rect 405 206 412 416
rect 395 199 412 206
rect 402 169 409 174
rect 395 167 409 169
rect 402 158 409 167
rect 402 120 409 128
<< ndiffusion >>
rect 136 275 157 297
rect 152 267 157 275
rect 164 267 197 297
rect 204 281 211 297
rect 227 281 238 297
rect 204 267 238 281
rect 245 267 279 297
rect 286 281 291 297
rect 286 267 307 281
rect 88 217 93 247
rect 100 217 157 247
rect 164 231 175 247
rect 164 217 191 231
rect 58 169 60 199
rect 67 169 72 199
rect 367 231 369 247
rect 351 217 369 231
rect 376 226 382 247
rect 376 217 398 226
rect 155 169 157 199
rect 164 169 197 199
rect 204 169 207 199
rect 271 169 279 199
rect 286 169 337 199
rect 344 169 348 199
rect 88 127 93 157
rect 100 141 105 157
rect 100 127 121 141
rect 236 141 238 157
rect 220 127 238 141
rect 245 127 279 157
rect 286 127 290 157
rect 399 128 402 158
rect 409 128 412 158
<< pdiffusion >>
rect 91 481 93 529
rect 100 481 102 529
rect 118 481 123 529
rect 130 503 148 529
rect 130 481 132 503
rect 57 419 60 464
rect 41 416 60 419
rect 67 437 88 464
rect 67 416 72 437
rect 262 481 279 529
rect 286 481 296 529
rect 312 481 337 529
rect 344 503 363 529
rect 344 481 347 503
rect 121 447 123 464
rect 105 416 123 447
rect 130 427 158 464
rect 174 427 176 464
rect 130 416 176 427
rect 183 427 196 464
rect 214 427 217 464
rect 183 416 217 427
rect 224 444 279 464
rect 224 427 226 444
rect 242 427 279 444
rect 224 416 279 427
rect 286 447 288 464
rect 286 416 299 447
rect 386 444 405 464
rect 75 370 93 396
rect 91 348 93 370
rect 100 348 103 396
rect 119 348 123 396
rect 130 348 132 396
rect 152 348 176 396
rect 183 390 217 396
rect 183 348 191 390
rect 209 348 217 390
rect 224 368 279 396
rect 224 348 226 368
rect 242 348 279 368
rect 286 390 305 396
rect 286 348 289 390
rect 402 416 405 444
rect 412 416 422 464
rect 350 390 369 396
rect 366 348 369 390
rect 376 370 394 396
rect 376 348 378 370
<< ntransistor >>
rect 157 267 164 297
rect 197 267 204 297
rect 238 267 245 297
rect 279 267 286 297
rect 93 217 100 247
rect 157 217 164 247
rect 60 169 67 199
rect 369 217 376 247
rect 157 169 164 199
rect 197 169 204 199
rect 279 169 286 199
rect 337 169 344 199
rect 93 127 100 157
rect 238 127 245 157
rect 279 127 286 157
rect 402 128 409 158
<< ptransistor >>
rect 93 481 100 529
rect 123 481 130 529
rect 60 416 67 464
rect 279 481 286 529
rect 337 481 344 529
rect 123 416 130 464
rect 176 416 183 464
rect 217 416 224 464
rect 279 416 286 464
rect 93 348 100 396
rect 123 348 130 396
rect 176 348 183 396
rect 217 348 224 396
rect 279 348 286 396
rect 405 416 412 464
rect 369 348 376 396
<< polycontact >>
rect 153 513 169 529
rect 208 480 224 496
rect 396 513 412 529
rect 360 421 376 437
rect 332 401 348 417
rect 176 322 192 338
rect 51 288 67 304
rect 89 288 105 304
rect 279 322 295 338
rect 281 210 297 226
rect 360 281 376 297
rect 229 169 245 199
rect 152 120 168 136
rect 193 120 210 137
rect 337 128 353 158
rect 386 169 402 199
<< ndiffcontact >>
rect 136 259 152 275
rect 211 281 227 297
rect 291 281 307 297
rect 72 217 88 247
rect 175 231 191 247
rect 42 169 58 199
rect 72 169 88 199
rect 351 231 367 247
rect 382 226 398 247
rect 139 169 155 199
rect 207 169 223 199
rect 255 169 271 199
rect 348 169 364 199
rect 72 127 88 157
rect 105 141 121 157
rect 220 141 236 157
rect 290 127 306 157
rect 383 128 399 158
rect 412 128 428 158
<< pdiffcontact >>
rect 75 481 91 529
rect 102 481 118 529
rect 132 481 148 503
rect 41 419 57 464
rect 72 416 88 437
rect 246 481 262 529
rect 296 481 312 529
rect 347 481 363 503
rect 105 447 121 464
rect 158 427 174 464
rect 196 427 214 464
rect 226 427 242 444
rect 288 447 304 464
rect 75 348 91 370
rect 103 348 119 396
rect 132 348 152 396
rect 191 348 209 390
rect 226 348 242 368
rect 289 348 305 390
rect 386 416 402 444
rect 350 348 366 390
rect 378 348 394 370
rect 422 415 438 464
<< psubstratetap >>
rect 246 89 263 106
<< nsubstratetap >>
rect 256 547 273 564
<< metal1 >>
rect 16 603 445 613
rect 16 579 335 589
rect 351 579 445 589
rect 16 564 445 566
rect 16 547 256 564
rect 273 547 445 564
rect 16 541 445 547
rect 41 464 57 541
rect 75 529 91 541
rect 118 519 153 529
rect 57 447 105 457
rect 132 457 142 481
rect 121 447 142 457
rect 158 480 208 490
rect 312 519 335 529
rect 350 519 396 529
rect 158 464 174 480
rect 246 464 262 481
rect 347 464 363 481
rect 422 464 438 541
rect 41 396 57 419
rect 88 427 158 437
rect 214 454 288 464
rect 304 454 422 464
rect 242 427 360 437
rect 132 401 306 411
rect 322 401 332 411
rect 386 411 402 416
rect 348 401 402 411
rect 132 396 152 401
rect 41 380 103 396
rect 422 390 438 415
rect 209 380 289 390
rect 305 380 350 390
rect 366 380 438 390
rect 75 338 91 348
rect 226 338 242 348
rect 378 338 394 348
rect 75 328 176 338
rect 192 328 242 338
rect 295 328 394 338
rect 30 291 51 301
rect 89 287 105 288
rect 115 297 227 303
rect 115 285 211 297
rect 115 247 126 285
rect 307 281 360 297
rect 152 259 428 269
rect 42 217 72 247
rect 88 237 126 247
rect 191 237 351 247
rect 88 217 271 219
rect 42 209 271 217
rect 382 221 398 226
rect 297 210 398 221
rect 42 199 58 209
rect 255 199 271 209
rect 88 169 139 199
rect 223 169 229 199
rect 364 169 386 199
rect 42 157 58 169
rect 412 158 428 259
rect 42 127 72 157
rect 121 147 220 157
rect 42 110 60 127
rect 151 120 152 136
rect 210 127 290 131
rect 353 128 383 158
rect 210 120 306 127
rect 30 106 445 110
rect 30 89 246 106
rect 263 89 445 106
rect 30 85 445 89
rect 30 61 89 71
rect 105 61 445 71
rect 30 38 445 48
rect 30 14 135 24
rect 151 14 445 24
<< m2contact >>
rect 335 576 351 592
rect 335 513 350 529
rect 306 401 322 417
rect 89 271 105 287
rect 135 120 151 136
rect 89 58 105 74
rect 135 10 151 26
<< metal2 >>
rect 308 417 320 625
rect 337 592 349 625
rect 337 529 349 576
rect 89 74 105 271
rect 135 26 151 120
rect 308 0 320 401
rect 337 0 349 513
<< labels >>
rlabel metal1 16 603 16 613 3 ScanReturn
rlabel metal1 16 579 16 589 3 Q
rlabel metal1 16 541 16 566 3 Vdd!
rlabel metal1 30 85 30 110 3 GND!
rlabel metal1 30 14 30 24 3 nRst
rlabel metal1 30 38 30 48 3 Test
rlabel metal1 30 61 30 71 3 Clk
rlabel metal1 30 291 30 301 3 D
rlabel metal2 337 0 349 0 1 Q
rlabel metal2 308 0 320 0 1 nQ
rlabel metal2 337 625 349 625 5 Q
rlabel metal2 308 625 320 625 5 nQ
<< end >>
