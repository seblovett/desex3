magic
tech c035u
timestamp 1386234512
<< nwell >>
rect 0 401 432 799
<< pwell >>
rect 0 0 432 401
<< polysilicon >>
rect 67 691 74 719
rect 97 691 104 719
rect 148 704 215 711
rect 34 610 41 621
rect 34 388 41 562
rect 67 486 74 643
rect 97 612 104 643
rect 150 612 157 623
rect 191 612 198 645
rect 208 624 215 704
rect 253 691 260 719
rect 311 691 318 719
rect 253 624 260 643
rect 208 617 260 624
rect 253 612 260 617
rect 97 486 104 564
rect 150 486 157 564
rect 191 486 198 564
rect 253 486 260 564
rect 311 532 318 643
rect 379 612 386 675
rect 34 220 41 372
rect 67 331 74 438
rect 97 402 104 438
rect 150 428 157 438
rect 166 412 178 419
rect 97 395 138 402
rect 131 358 138 395
rect 171 358 178 412
rect 191 410 198 438
rect 253 428 260 438
rect 191 403 219 410
rect 212 358 219 403
rect 253 358 260 412
rect 67 288 74 315
rect 131 288 138 328
rect 34 182 41 190
rect 67 161 74 258
rect 131 220 138 258
rect 171 220 178 328
rect 212 220 219 328
rect 253 255 260 328
rect 253 248 267 255
rect 253 225 267 232
rect 253 220 260 225
rect 311 220 318 516
rect 343 486 350 539
rect 343 358 350 438
rect 343 288 350 328
rect 67 110 74 131
rect 131 127 138 190
rect 171 128 178 190
rect 212 161 219 190
rect 253 161 260 190
rect 311 180 318 190
rect 311 142 318 150
rect 343 142 350 258
rect 379 227 386 564
rect 369 220 386 227
rect 376 190 383 195
rect 369 188 383 190
rect 376 180 383 188
rect 376 142 383 150
rect 212 120 219 131
rect 253 120 260 131
<< ndiffusion >>
rect 126 328 131 358
rect 138 328 171 358
rect 178 328 185 358
rect 201 328 212 358
rect 219 328 253 358
rect 260 328 265 358
rect 62 258 67 288
rect 74 258 131 288
rect 138 258 149 288
rect 32 190 34 220
rect 41 190 46 220
rect 341 258 343 288
rect 350 258 356 288
rect 129 190 131 220
rect 138 190 171 220
rect 178 190 181 220
rect 245 190 253 220
rect 260 190 311 220
rect 318 190 322 220
rect 62 131 67 161
rect 74 131 79 161
rect 210 131 212 161
rect 219 131 253 161
rect 260 131 264 161
rect 373 150 376 180
rect 383 150 386 180
<< pdiffusion >>
rect 65 643 67 691
rect 74 643 76 691
rect 92 643 97 691
rect 104 643 106 691
rect 31 562 34 610
rect 41 562 46 610
rect 236 643 253 691
rect 260 643 270 691
rect 286 643 311 691
rect 318 643 321 691
rect 95 564 97 612
rect 104 564 132 612
rect 148 564 150 612
rect 157 564 167 612
rect 183 564 191 612
rect 198 564 200 612
rect 216 564 253 612
rect 260 564 262 612
rect 376 564 379 612
rect 386 564 396 612
rect 65 438 67 486
rect 74 438 77 486
rect 93 438 97 486
rect 104 438 106 486
rect 126 438 150 486
rect 157 438 165 486
rect 183 438 191 486
rect 198 438 200 486
rect 216 438 253 486
rect 260 438 263 486
rect 340 438 343 486
rect 350 438 356 486
<< pohmic >>
rect 0 76 10 86
rect 26 76 38 86
rect 54 76 66 86
rect 82 76 94 86
rect 110 76 122 86
rect 138 76 150 86
rect 166 76 178 86
rect 194 76 206 86
rect 222 76 234 86
rect 251 76 263 86
rect 279 76 291 86
rect 307 76 319 86
rect 335 76 347 86
rect 364 76 376 86
rect 393 76 405 86
rect 422 76 432 86
<< nohmic >>
rect 0 736 10 746
rect 26 736 38 746
rect 54 736 66 746
rect 82 736 94 746
rect 110 736 122 746
rect 138 736 150 746
rect 166 736 178 746
rect 194 736 206 746
rect 222 736 234 746
rect 250 736 262 746
rect 278 736 290 746
rect 306 736 318 746
rect 334 736 346 746
rect 362 736 374 746
rect 390 736 402 746
rect 418 736 432 746
<< ntransistor >>
rect 131 328 138 358
rect 171 328 178 358
rect 212 328 219 358
rect 253 328 260 358
rect 67 258 74 288
rect 131 258 138 288
rect 34 190 41 220
rect 343 258 350 288
rect 131 190 138 220
rect 171 190 178 220
rect 253 190 260 220
rect 311 190 318 220
rect 67 131 74 161
rect 212 131 219 161
rect 253 131 260 161
rect 376 150 383 180
<< ptransistor >>
rect 67 643 74 691
rect 97 643 104 691
rect 34 562 41 610
rect 253 643 260 691
rect 311 643 318 691
rect 97 564 104 612
rect 150 564 157 612
rect 191 564 198 612
rect 253 564 260 612
rect 379 564 386 612
rect 67 438 74 486
rect 97 438 104 486
rect 150 438 157 486
rect 191 438 198 486
rect 253 438 260 486
rect 343 438 350 486
<< polycontact >>
rect 132 695 148 711
rect 182 645 198 661
rect 370 675 386 691
rect 334 539 350 555
rect 306 516 322 532
rect 25 372 41 388
rect 150 412 166 428
rect 253 412 269 428
rect 63 315 79 331
rect 255 232 271 248
rect 334 328 350 358
rect 203 190 219 220
rect 311 150 327 180
rect 360 190 376 220
rect 126 111 142 127
rect 167 111 184 128
<< ndiffcontact >>
rect 110 328 126 358
rect 185 328 201 358
rect 265 328 281 358
rect 46 258 62 288
rect 149 258 165 288
rect 16 190 32 220
rect 46 190 62 220
rect 325 258 341 288
rect 356 258 372 288
rect 113 190 129 220
rect 181 190 197 220
rect 229 190 245 220
rect 322 190 338 220
rect 46 131 62 161
rect 79 131 95 161
rect 194 131 210 161
rect 264 131 280 161
rect 357 150 373 180
rect 386 150 402 180
<< pdiffcontact >>
rect 49 643 65 691
rect 76 643 92 691
rect 106 643 122 691
rect 15 562 31 610
rect 46 562 62 610
rect 220 643 236 691
rect 270 643 286 691
rect 321 643 337 691
rect 79 564 95 612
rect 132 564 148 612
rect 167 564 183 612
rect 200 564 216 612
rect 262 564 278 612
rect 360 564 376 612
rect 396 564 412 612
rect 49 438 65 486
rect 77 438 93 486
rect 106 438 126 486
rect 165 438 183 486
rect 200 438 216 486
rect 263 438 279 486
rect 324 438 340 486
rect 356 438 373 486
<< psubstratetap >>
rect 10 76 26 92
rect 38 76 54 92
rect 66 76 82 92
rect 94 76 110 92
rect 122 76 138 92
rect 150 76 166 92
rect 178 76 194 92
rect 206 76 222 92
rect 234 76 251 92
rect 263 76 279 92
rect 291 76 307 92
rect 319 76 335 92
rect 347 76 364 92
rect 376 76 393 92
rect 405 76 422 92
<< nsubstratetap >>
rect 10 730 26 746
rect 38 730 54 746
rect 66 730 82 746
rect 94 730 110 746
rect 122 730 138 746
rect 150 730 166 746
rect 178 730 194 746
rect 206 730 222 746
rect 234 730 250 746
rect 262 730 278 746
rect 290 730 306 746
rect 318 730 334 746
rect 346 730 362 746
rect 374 730 390 746
rect 402 730 418 746
<< metal1 >>
rect 0 782 432 792
rect 0 759 314 769
rect 330 759 432 769
rect 0 730 10 746
rect 26 730 38 746
rect 54 730 66 746
rect 82 730 94 746
rect 110 730 122 746
rect 138 730 150 746
rect 166 730 178 746
rect 194 730 206 746
rect 222 730 234 746
rect 250 730 262 746
rect 278 730 290 746
rect 306 730 318 746
rect 334 730 346 746
rect 362 730 374 746
rect 390 730 402 746
rect 418 730 432 746
rect 0 721 432 730
rect 15 634 31 721
rect 49 691 65 721
rect 76 701 132 711
rect 76 691 92 701
rect 270 701 370 711
rect 270 691 286 701
rect 370 691 386 695
rect 15 633 32 634
rect 106 633 122 643
rect 15 621 122 633
rect 132 645 182 655
rect 15 610 31 621
rect 79 612 95 621
rect 15 511 31 562
rect 132 612 148 645
rect 220 633 236 643
rect 321 633 337 643
rect 396 633 412 721
rect 167 623 412 633
rect 167 612 183 623
rect 262 612 278 623
rect 396 612 412 623
rect 46 549 62 562
rect 132 549 148 564
rect 46 539 148 549
rect 200 554 216 564
rect 200 544 334 554
rect 106 516 266 526
rect 282 516 306 526
rect 360 526 376 564
rect 322 516 376 526
rect 15 501 93 511
rect 77 486 93 501
rect 106 486 126 516
rect 396 506 412 564
rect 165 496 279 506
rect 165 486 183 496
rect 263 486 279 496
rect 324 496 412 506
rect 324 486 340 496
rect 279 438 324 486
rect 49 428 65 438
rect 200 428 216 438
rect 356 428 373 438
rect 49 418 150 428
rect 166 418 216 428
rect 269 418 373 428
rect 64 390 201 402
rect 0 375 25 385
rect 64 353 77 390
rect 185 358 201 390
rect 16 341 77 353
rect 16 288 32 341
rect 63 314 79 315
rect 281 328 334 358
rect 110 318 126 328
rect 110 308 402 318
rect 16 258 46 288
rect 165 278 325 288
rect 16 220 32 258
rect 46 247 62 258
rect 356 248 372 258
rect 46 235 245 247
rect 229 220 245 235
rect 271 232 372 248
rect 62 190 113 220
rect 197 190 203 220
rect 338 190 360 220
rect 16 161 32 190
rect 386 180 402 308
rect 16 131 46 161
rect 95 151 194 161
rect 327 150 357 180
rect 16 101 34 131
rect 125 111 126 127
rect 264 121 280 131
rect 184 111 280 121
rect 0 92 432 101
rect 0 76 10 92
rect 26 76 38 92
rect 54 76 66 92
rect 82 76 94 92
rect 110 76 122 92
rect 138 76 150 92
rect 166 76 178 92
rect 194 76 206 92
rect 222 76 234 92
rect 251 76 263 92
rect 279 76 291 92
rect 307 76 319 92
rect 335 76 347 92
rect 364 76 376 92
rect 393 76 405 92
rect 422 76 432 92
rect 0 53 63 63
rect 79 53 432 63
rect 0 30 432 40
rect 0 7 109 17
rect 125 7 432 17
<< m2contact >>
rect 314 756 330 772
rect 370 695 386 711
rect 266 516 282 532
rect 63 298 79 314
rect 109 111 125 127
rect 63 50 79 66
rect 109 4 125 20
<< metal2 >>
rect 268 532 280 799
rect 316 772 328 799
rect 316 711 328 756
rect 316 695 370 711
rect 63 66 79 298
rect 109 20 125 111
rect 268 0 280 516
rect 316 0 328 695
<< labels >>
rlabel metal2 268 799 280 799 5 nQ
rlabel metal2 268 0 280 0 1 nQ
rlabel metal2 316 799 328 799 5 Q
rlabel metal2 316 0 328 0 1 Q
rlabel metal1 0 375 0 385 3 D
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 759 0 769 3 Q
rlabel metal1 0 7 0 17 1 nReset
rlabel metal1 0 53 0 63 1 Clock
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 432 782 432 792 7 ScanReturn
rlabel metal1 432 759 432 769 7 Q
rlabel metal1 432 76 432 101 7 GND!
rlabel metal1 432 53 432 63 7 Clock
rlabel metal1 432 30 432 40 7 Test
rlabel metal1 432 7 432 17 7 nReset
rlabel metal1 432 721 432 746 7 Vdd!
<< end >>
