magic
tech c035u
timestamp 1384967361
<< nwell >>
rect 0 219 140 308
<< polysilicon >>
rect 28 274 35 282
rect 55 274 62 282
rect 82 274 89 282
rect 109 274 116 282
rect 28 94 35 226
rect 55 156 62 226
rect 61 140 62 156
rect 28 68 35 78
rect 55 68 62 140
rect 82 113 89 226
rect 109 154 116 226
rect 115 138 116 154
rect 108 124 116 138
rect 88 97 89 113
rect 81 83 89 97
rect 82 68 89 83
rect 109 68 116 124
rect 28 30 35 38
rect 55 30 62 38
rect 82 30 89 38
rect 109 30 116 38
<< ndiffusion >>
rect 26 38 28 68
rect 35 38 55 68
rect 62 38 82 68
rect 89 38 109 68
rect 116 38 118 68
<< pdiffusion >>
rect 26 226 28 274
rect 35 226 37 274
rect 53 226 55 274
rect 62 226 64 274
rect 80 226 82 274
rect 89 226 91 274
rect 107 226 109 274
rect 116 226 118 274
<< pohmic >>
rect 0 7 6 14
rect 22 7 34 14
rect 50 7 62 14
rect 78 7 90 14
rect 106 7 118 14
rect 134 7 140 14
rect 0 4 140 7
<< nohmic >>
rect 0 305 140 308
rect 0 298 6 305
rect 22 298 34 305
rect 50 298 62 305
rect 78 298 90 305
rect 106 298 118 305
rect 134 298 140 305
<< ntransistor >>
rect 28 38 35 68
rect 55 38 62 68
rect 82 38 89 68
rect 109 38 116 68
<< ptransistor >>
rect 28 226 35 274
rect 55 226 62 274
rect 82 226 89 274
rect 109 226 116 274
<< polycontact >>
rect 45 140 61 156
rect 24 78 40 94
rect 99 138 115 154
rect 72 97 88 113
<< ndiffcontact >>
rect 10 38 26 68
rect 118 38 134 68
<< pdiffcontact >>
rect 10 226 26 274
rect 37 226 53 274
rect 64 226 80 274
rect 91 226 107 274
rect 118 226 134 274
<< psubstratetap >>
rect 6 7 22 23
rect 34 7 50 23
rect 62 7 78 23
rect 90 7 106 23
rect 118 7 134 23
<< nsubstratetap >>
rect 6 289 22 305
rect 34 289 50 305
rect 62 289 78 305
rect 90 289 106 305
rect 118 289 134 305
<< metal1 >>
rect 0 305 140 308
rect 0 289 6 305
rect 22 289 34 305
rect 50 289 62 305
rect 78 289 90 305
rect 106 289 118 305
rect 134 289 140 305
rect 0 284 140 289
rect 10 274 26 284
rect 64 274 80 284
rect 118 274 134 284
rect 43 176 53 226
rect 97 176 107 226
rect 43 166 121 176
rect 125 68 135 164
rect 134 38 135 68
rect 10 28 26 38
rect 0 23 140 28
rect 0 7 6 23
rect 22 7 34 23
rect 50 7 62 23
rect 78 7 90 23
rect 106 7 118 23
rect 134 7 140 23
rect 0 4 140 7
<< m2contact >>
rect 121 164 135 178
rect 46 126 60 140
rect 96 124 110 138
rect 24 94 38 108
rect 72 83 86 97
<< metal2 >>
rect 24 274 36 312
rect 24 226 37 274
rect 24 108 36 226
rect 48 156 60 312
rect 48 140 61 156
rect 24 78 38 94
rect 24 23 36 78
rect 23 7 36 23
rect 24 0 36 7
rect 48 0 60 126
rect 72 97 84 312
rect 96 274 108 312
rect 96 226 109 274
rect 96 138 108 226
rect 120 178 132 311
rect 120 164 121 178
rect 72 0 84 83
rect 96 0 108 124
rect 120 68 132 164
rect 120 38 134 68
rect 120 0 132 38
<< labels >>
rlabel metal1 0 284 0 308 3 Vdd!
rlabel metal2 24 312 36 312 5 A
rlabel metal2 48 312 60 312 5 B
rlabel metal2 48 0 60 0 1 B
rlabel metal2 24 0 36 0 1 A
rlabel metal1 0 4 0 28 3 GND!
rlabel metal2 72 312 84 312 5 C
rlabel metal2 72 0 84 0 1 C
rlabel metal2 96 0 108 0 1 D
rlabel metal2 96 312 108 312 5 D
rlabel metal2 120 0 132 0 1 Y
rlabel metal1 140 4 140 28 7 GND!
rlabel metal1 140 284 140 308 7 Vdd!
<< end >>
