magic
tech c035u
timestamp 1386265531
<< nwell >>
rect 0 427 672 825
<< pwell >>
rect 0 26 672 427
<< polysilicon >>
rect 275 656 282 664
rect 302 656 309 664
rect 333 656 340 664
rect 275 531 282 608
rect 302 572 309 608
rect 333 598 340 608
rect 395 607 404 614
rect 302 556 304 572
rect 302 531 309 556
rect 55 495 62 503
rect 175 495 182 503
rect 55 417 62 447
rect 175 417 182 447
rect 275 432 282 483
rect 273 423 282 432
rect 60 401 62 417
rect 180 401 182 417
rect 278 407 282 423
rect 55 366 62 401
rect 175 366 182 401
rect 275 392 282 407
rect 302 392 309 483
rect 333 392 340 582
rect 367 531 374 539
rect 397 531 404 607
rect 487 495 494 503
rect 607 495 614 503
rect 367 473 374 483
rect 55 328 62 336
rect 175 328 182 336
rect 275 319 282 362
rect 302 319 309 362
rect 333 319 340 371
rect 367 361 374 457
rect 397 361 404 483
rect 487 417 494 447
rect 607 417 614 447
rect 492 401 494 417
rect 612 401 614 417
rect 487 366 494 401
rect 607 366 614 401
rect 367 323 374 331
rect 397 313 404 331
rect 487 328 494 336
rect 607 328 614 336
rect 393 306 404 313
rect 275 281 282 289
rect 302 281 309 289
rect 333 281 340 289
<< ndiffusion >>
rect 53 336 55 366
rect 62 336 64 366
rect 173 336 175 366
rect 182 336 184 366
rect 272 362 275 392
rect 282 362 302 392
rect 309 362 311 392
rect 365 331 367 361
rect 374 331 378 361
rect 394 331 397 361
rect 404 331 406 361
rect 485 336 487 366
rect 494 336 496 366
rect 605 336 607 366
rect 614 336 616 366
rect 272 289 275 319
rect 282 289 284 319
rect 300 289 302 319
rect 309 289 311 319
rect 327 289 333 319
rect 340 289 342 319
<< pdiffusion >>
rect 273 608 275 656
rect 282 608 284 656
rect 300 608 302 656
rect 309 608 311 656
rect 327 608 333 656
rect 340 608 342 656
rect 53 447 55 495
rect 62 447 64 495
rect 173 447 175 495
rect 182 447 184 495
rect 273 483 275 531
rect 282 483 302 531
rect 309 483 312 531
rect 364 483 367 531
rect 374 483 397 531
rect 404 483 406 531
rect 485 447 487 495
rect 494 447 496 495
rect 605 447 607 495
rect 614 447 616 495
<< pohmic >>
rect 0 102 6 112
rect 22 102 34 112
rect 50 102 62 112
rect 78 102 90 112
rect 106 102 126 112
rect 142 102 154 112
rect 170 102 182 112
rect 198 102 210 112
rect 226 102 251 112
rect 267 102 279 112
rect 295 102 307 112
rect 323 102 335 112
rect 351 102 363 112
rect 379 102 391 112
rect 407 102 438 112
rect 454 102 466 112
rect 482 102 494 112
rect 510 102 522 112
rect 538 102 558 112
rect 574 102 586 112
rect 602 102 614 112
rect 630 102 642 112
rect 658 102 672 112
<< nohmic >>
rect 0 762 6 772
rect 22 762 34 772
rect 50 762 62 772
rect 78 762 90 772
rect 106 762 126 772
rect 142 762 154 772
rect 170 762 182 772
rect 198 762 210 772
rect 226 762 251 772
rect 267 762 279 772
rect 295 762 307 772
rect 323 762 335 772
rect 351 762 363 772
rect 379 762 391 772
rect 407 762 438 772
rect 454 762 466 772
rect 482 762 494 772
rect 510 762 522 772
rect 538 762 558 772
rect 574 762 586 772
rect 602 762 614 772
rect 630 762 642 772
rect 658 762 672 772
<< ntransistor >>
rect 55 336 62 366
rect 175 336 182 366
rect 275 362 282 392
rect 302 362 309 392
rect 367 331 374 361
rect 397 331 404 361
rect 487 336 494 366
rect 607 336 614 366
rect 275 289 282 319
rect 302 289 309 319
rect 333 289 340 319
<< ptransistor >>
rect 275 608 282 656
rect 302 608 309 656
rect 333 608 340 656
rect 55 447 62 495
rect 175 447 182 495
rect 275 483 282 531
rect 302 483 309 531
rect 367 483 374 531
rect 397 483 404 531
rect 487 447 494 495
rect 607 447 614 495
<< polycontact >>
rect 379 607 395 623
rect 325 582 341 598
rect 304 556 320 572
rect 44 401 60 417
rect 164 401 180 417
rect 262 407 278 423
rect 358 457 374 473
rect 333 371 349 392
rect 476 401 492 417
rect 596 401 612 417
rect 377 289 393 313
<< ndiffcontact >>
rect 37 336 53 366
rect 64 336 80 366
rect 157 336 173 366
rect 184 336 200 366
rect 256 362 272 392
rect 311 362 327 392
rect 349 331 365 361
rect 378 331 394 361
rect 406 331 422 361
rect 469 336 485 366
rect 496 336 512 366
rect 589 336 605 366
rect 616 336 632 366
rect 256 289 272 319
rect 284 289 300 319
rect 311 289 327 319
rect 342 289 358 319
<< pdiffcontact >>
rect 257 608 273 656
rect 284 608 300 656
rect 311 608 327 656
rect 342 608 358 656
rect 37 447 53 495
rect 64 447 80 495
rect 157 447 173 495
rect 184 447 200 495
rect 257 483 273 531
rect 312 483 328 531
rect 348 483 364 531
rect 406 483 422 531
rect 469 447 485 495
rect 496 447 512 495
rect 589 447 605 495
rect 616 447 632 495
<< psubstratetap >>
rect 37 307 53 323
rect 157 307 173 323
rect 469 307 485 323
rect 589 307 605 323
rect 406 270 422 286
rect 406 242 422 258
rect 406 214 422 230
rect 406 186 422 202
rect 406 158 422 174
rect 406 130 422 146
rect 6 102 22 118
rect 34 102 50 118
rect 62 102 78 118
rect 90 102 106 118
rect 126 102 142 118
rect 154 102 170 118
rect 182 102 198 118
rect 210 102 226 118
rect 251 102 267 118
rect 279 102 295 118
rect 307 102 323 118
rect 335 102 351 118
rect 363 102 379 118
rect 391 102 407 118
rect 438 102 454 118
rect 466 102 482 118
rect 494 102 510 118
rect 522 102 538 118
rect 558 102 574 118
rect 586 102 602 118
rect 614 102 630 118
rect 642 102 658 118
<< nsubstratetap >>
rect 6 756 22 772
rect 34 756 50 772
rect 62 756 78 772
rect 90 756 106 772
rect 126 756 142 772
rect 154 756 170 772
rect 182 756 198 772
rect 210 756 226 772
rect 251 756 267 772
rect 279 756 295 772
rect 307 756 323 772
rect 335 756 351 772
rect 363 756 379 772
rect 391 756 407 772
rect 438 756 454 772
rect 466 756 482 772
rect 494 756 510 772
rect 522 756 538 772
rect 558 756 574 772
rect 586 756 602 772
rect 614 756 630 772
rect 642 756 658 772
<< metal1 >>
rect 397 865 455 875
rect 469 865 575 875
rect 205 844 263 854
rect 0 808 672 818
rect 0 785 672 795
rect 0 756 6 772
rect 22 756 34 772
rect 50 756 62 772
rect 78 756 90 772
rect 106 756 126 772
rect 142 756 154 772
rect 170 756 182 772
rect 198 756 210 772
rect 226 756 251 772
rect 267 756 279 772
rect 295 756 307 772
rect 323 756 335 772
rect 351 756 363 772
rect 379 756 391 772
rect 407 756 438 772
rect 454 756 466 772
rect 482 756 494 772
rect 510 756 522 772
rect 538 756 558 772
rect 574 756 586 772
rect 602 756 614 772
rect 630 756 642 772
rect 658 756 672 772
rect 0 747 672 756
rect 37 495 53 747
rect 157 495 173 747
rect 257 656 273 747
rect 311 656 327 747
rect 358 608 379 622
rect 257 531 273 608
rect 287 595 297 608
rect 287 585 325 595
rect 406 531 423 747
rect 364 483 394 493
rect 422 483 423 531
rect 469 495 485 747
rect 589 495 605 747
rect 312 471 328 483
rect 70 415 80 447
rect 190 415 200 447
rect 290 459 358 471
rect 262 423 278 424
rect 70 366 80 401
rect 190 366 200 401
rect 37 323 53 336
rect 37 127 53 307
rect 157 323 173 336
rect 157 127 173 307
rect 256 319 272 362
rect 290 319 300 459
rect 384 420 394 483
rect 327 371 333 392
rect 384 361 394 404
rect 502 415 512 447
rect 622 415 632 447
rect 502 366 512 401
rect 622 366 632 401
rect 311 331 349 350
rect 311 319 327 331
rect 358 289 377 313
rect 256 127 272 289
rect 311 127 327 289
rect 406 286 422 331
rect 406 258 422 270
rect 406 230 422 242
rect 406 202 422 214
rect 406 174 422 186
rect 406 146 422 158
rect 406 127 422 130
rect 469 323 485 336
rect 469 127 485 307
rect 589 323 605 336
rect 589 127 605 307
rect 0 118 672 127
rect 0 102 6 118
rect 22 102 34 118
rect 50 102 62 118
rect 78 102 90 118
rect 106 102 126 118
rect 142 102 154 118
rect 170 102 182 118
rect 198 102 210 118
rect 226 102 251 118
rect 267 102 279 118
rect 295 102 307 118
rect 323 102 335 118
rect 351 102 363 118
rect 379 102 391 118
rect 407 102 438 118
rect 454 102 466 118
rect 482 102 494 118
rect 510 102 522 118
rect 538 102 558 118
rect 574 102 586 118
rect 602 102 614 118
rect 630 102 642 118
rect 658 102 672 118
rect 0 79 672 89
rect 0 56 672 66
rect 0 33 672 43
rect 85 2 287 12
<< m2contact >>
rect 383 863 397 877
rect 455 863 469 877
rect 575 863 589 877
rect 191 842 205 856
rect 263 842 277 856
rect 288 556 304 572
rect 30 402 44 416
rect 70 401 84 415
rect 150 402 164 416
rect 262 424 278 440
rect 190 401 204 415
rect 381 404 397 420
rect 462 402 476 416
rect 502 401 516 415
rect 582 402 596 416
rect 622 401 636 415
rect 71 0 85 14
rect 287 0 301 14
<< metal2 >>
rect 24 416 36 911
rect 24 402 30 416
rect 72 415 84 825
rect 24 26 36 402
rect 72 14 84 401
rect 144 416 156 911
rect 264 856 276 911
rect 144 402 150 416
rect 192 415 204 842
rect 264 440 276 842
rect 288 572 300 911
rect 384 877 396 911
rect 304 558 305 572
rect 262 423 276 424
rect 144 26 156 402
rect 192 26 204 401
rect 264 26 276 423
rect 288 14 300 556
rect 384 420 396 863
rect 456 416 468 863
rect 384 26 396 404
rect 456 402 462 416
rect 504 415 516 825
rect 456 26 468 402
rect 504 26 516 401
rect 576 416 588 863
rect 576 402 582 416
rect 624 415 636 825
rect 576 26 588 402
rect 624 26 636 401
<< labels >>
rlabel metal1 672 747 672 772 7 Vdd!
rlabel metal1 672 785 672 795 7 Scan
rlabel metal1 672 808 672 818 6 ScanReturn
rlabel metal1 672 33 672 43 8 nReset
rlabel metal1 672 56 672 66 7 Test
rlabel metal1 672 79 672 89 7 Clock
rlabel metal1 672 102 672 127 7 GND!
rlabel metal2 24 911 36 911 5 nB
rlabel metal2 144 911 156 911 5 nA
rlabel metal2 264 911 276 911 5 A
rlabel metal2 288 911 300 911 5 B
rlabel metal2 384 911 396 911 5 Y
<< end >>
