magic
tech c035u
timestamp 1385123640
<< nwell >>
rect 0 460 192 659
<< polysilicon >>
rect 29 604 36 612
rect 59 604 66 612
rect 92 604 99 612
rect 119 604 126 612
rect 150 604 157 612
rect 29 525 36 556
rect 59 512 66 556
rect 92 509 99 556
rect 29 270 36 477
rect 59 270 66 496
rect 119 504 126 556
rect 150 546 157 556
rect 153 530 157 546
rect 92 270 99 493
rect 119 270 126 488
rect 150 316 157 530
rect 152 300 157 316
rect 29 209 36 244
rect 59 205 66 244
rect 92 236 99 244
rect 119 236 126 244
rect 150 209 157 300
rect 29 173 36 183
rect 150 175 157 183
rect 29 157 37 173
<< ndiffusion >>
rect 27 244 29 270
rect 36 244 38 270
rect 54 244 59 270
rect 66 244 92 270
rect 99 244 101 270
rect 117 244 119 270
rect 126 244 128 270
rect 27 183 29 209
rect 36 183 38 209
rect 148 183 150 209
rect 157 183 159 209
<< pdiffusion >>
rect 27 556 29 604
rect 36 556 38 604
rect 54 556 59 604
rect 66 556 68 604
rect 84 556 92 604
rect 99 556 101 604
rect 117 556 119 604
rect 126 556 129 604
rect 145 556 150 604
rect 157 556 160 604
rect 27 477 29 525
rect 36 477 38 525
<< pohmic >>
rect 0 2 6 9
rect 22 2 34 9
rect 50 2 62 9
rect 78 2 90 9
rect 106 2 118 9
rect 134 2 146 9
rect 162 2 192 9
rect 0 -1 192 2
<< nohmic >>
rect 0 656 192 659
rect 0 649 8 656
rect 24 649 36 656
rect 52 649 64 656
rect 80 649 92 656
rect 108 649 120 656
rect 136 649 148 656
rect 164 649 192 656
<< ntransistor >>
rect 29 244 36 270
rect 59 244 66 270
rect 92 244 99 270
rect 119 244 126 270
rect 29 183 36 209
rect 150 183 157 209
<< ptransistor >>
rect 29 556 36 604
rect 59 556 66 604
rect 92 556 99 604
rect 119 556 126 604
rect 150 556 157 604
rect 29 477 36 525
<< polycontact >>
rect 59 496 75 512
rect 88 493 104 509
rect 137 530 153 546
rect 117 488 133 504
rect 136 300 152 316
rect 59 189 75 205
rect 37 157 53 173
<< ndiffcontact >>
rect 11 244 27 270
rect 38 244 54 270
rect 101 244 117 270
rect 128 244 144 270
rect 11 183 27 209
rect 38 183 54 209
rect 132 183 148 209
rect 159 183 175 209
<< pdiffcontact >>
rect 11 556 27 604
rect 38 556 54 604
rect 68 556 84 604
rect 101 556 117 604
rect 129 556 145 604
rect 160 556 176 604
rect 11 477 27 525
rect 38 477 54 525
<< psubstratetap >>
rect 6 2 22 18
rect 34 2 50 18
rect 62 2 78 18
rect 90 2 106 18
rect 118 2 134 18
rect 146 2 162 18
<< nsubstratetap >>
rect 8 640 24 656
rect 36 640 52 656
rect 64 640 80 656
rect 92 640 108 656
rect 120 640 136 656
rect 148 640 164 656
<< metal1 >>
rect 0 695 192 705
rect 0 672 120 682
rect 0 656 192 659
rect 0 640 8 656
rect 24 640 36 656
rect 52 640 64 656
rect 80 640 92 656
rect 108 640 120 656
rect 136 640 148 656
rect 164 640 192 656
rect 0 634 192 640
rect 11 604 27 634
rect 41 614 114 624
rect 41 604 51 614
rect 104 604 114 614
rect 129 604 145 634
rect 11 525 27 556
rect 71 542 81 556
rect 71 532 137 542
rect 54 496 59 512
rect 163 385 173 556
rect 163 375 192 385
rect 41 303 136 313
rect 41 270 51 303
rect 73 280 141 290
rect 14 234 24 244
rect 73 234 83 280
rect 131 270 141 280
rect 14 224 83 234
rect 54 189 59 205
rect 11 24 27 183
rect 101 24 117 244
rect 163 209 173 375
rect 132 24 148 183
rect 0 18 192 24
rect 0 2 6 18
rect 22 2 34 18
rect 50 2 62 18
rect 78 2 90 18
rect 106 2 118 18
rect 134 2 146 18
rect 162 2 192 18
rect 0 -1 192 2
rect 0 -24 192 -14
rect 0 -47 39 -37
rect 53 -47 192 -37
rect 0 -70 192 -60
<< m2contact >>
rect 120 670 134 684
rect 119 504 133 518
rect 89 479 103 493
rect 39 143 53 157
rect 39 -49 53 -35
<< metal2 >>
rect 97 493 109 709
rect 121 518 133 670
rect 103 479 109 493
rect 40 -35 52 143
rect 97 -74 109 479
<< labels >>
rlabel metal1 0 -1 0 24 1 GND!
rlabel metal1 0 -70 0 -60 2 nReset
rlabel metal1 0 -47 0 -37 3 Test
rlabel metal1 0 -24 0 -14 3 Clock
rlabel metal1 0 634 0 659 3 Vdd!
rlabel metal1 0 672 0 682 3 Scan
rlabel metal1 0 695 0 705 4 ScanReturn
rlabel metal2 97 -74 109 -74 1 D
rlabel metal2 97 709 109 709 5 D
rlabel metal1 192 375 192 385 7 M
rlabel metal1 192 -1 192 24 7 GND!
rlabel metal1 192 -70 192 -60 8 nReset
rlabel metal1 192 -47 192 -37 7 Test
rlabel metal1 192 -24 192 -14 7 Clock
rlabel metal1 192 634 192 659 7 Vdd!
rlabel metal1 192 695 192 705 6 ScanReturn
<< end >>
