magic
tech c035u
timestamp 1385074831
<< nwell >>
rect 3 483 340 728
rect 3 482 327 483
rect 35 390 327 482
rect 88 389 134 390
<< polysilicon >>
rect 221 680 228 688
rect 248 680 255 688
rect 275 680 282 688
rect 302 680 309 688
rect 163 602 170 610
rect 190 602 197 610
rect 53 448 60 576
rect 108 547 115 555
rect 53 376 60 390
rect 108 376 115 390
rect 163 377 170 390
rect 58 360 60 376
rect 113 360 115 376
rect 168 373 170 377
rect 190 373 197 390
rect 221 377 228 390
rect 168 366 197 373
rect 168 361 170 366
rect 226 373 228 377
rect 248 373 255 390
rect 275 373 282 390
rect 302 373 309 390
rect 226 366 309 373
rect 226 361 228 366
rect 53 350 60 360
rect 108 350 115 360
rect 163 350 170 361
rect 221 350 228 361
rect 248 350 255 366
rect 53 322 60 330
rect 108 288 115 296
rect 163 196 170 204
rect 221 142 228 150
rect 248 142 255 150
<< ndiffusion >>
rect 51 330 53 350
rect 60 330 62 350
rect 106 296 108 350
rect 115 296 117 350
rect 161 204 163 350
rect 170 204 172 350
rect 219 150 221 350
rect 228 150 230 350
rect 246 150 248 350
rect 255 150 257 350
<< pdiffusion >>
rect 51 390 53 448
rect 60 390 62 448
rect 106 390 108 547
rect 115 390 117 547
rect 161 390 163 602
rect 170 390 172 602
rect 188 390 190 602
rect 197 390 199 602
rect 219 390 221 680
rect 228 390 230 680
rect 246 390 248 680
rect 255 390 257 680
rect 273 390 275 680
rect 282 390 284 680
rect 300 390 302 680
rect 309 390 311 680
<< pohmic >>
rect 3 70 9 80
rect 25 70 37 80
rect 53 70 65 80
rect 81 70 93 80
rect 109 70 121 80
rect 137 70 149 80
rect 165 70 177 80
rect 193 70 205 80
rect 221 70 233 80
rect 250 70 262 80
rect 278 70 290 80
rect 306 70 318 80
rect 334 70 340 80
<< nohmic >>
rect 3 718 9 728
rect 25 718 37 728
rect 53 718 65 728
rect 81 718 93 728
rect 109 718 121 728
rect 137 718 149 728
rect 165 718 177 728
rect 193 718 205 728
rect 221 718 233 728
rect 250 718 262 728
rect 278 718 290 728
rect 306 718 318 728
rect 334 718 340 728
<< ntransistor >>
rect 53 330 60 350
rect 108 296 115 350
rect 163 204 170 350
rect 221 150 228 350
rect 248 150 255 350
<< ptransistor >>
rect 53 390 60 448
rect 108 390 115 547
rect 163 390 170 602
rect 190 390 197 602
rect 221 390 228 680
rect 248 390 255 680
rect 275 390 282 680
rect 302 390 309 680
<< polycontact >>
rect 42 360 58 376
rect 97 360 113 376
rect 152 361 168 377
rect 210 361 226 377
<< ndiffcontact >>
rect 35 330 51 350
rect 62 330 78 350
rect 90 296 106 350
rect 117 296 133 350
rect 145 204 161 350
rect 172 204 188 350
rect 203 150 219 350
rect 230 150 246 350
rect 257 150 273 350
<< pdiffcontact >>
rect 202 602 219 680
rect 35 390 51 448
rect 62 390 78 448
rect 90 390 106 547
rect 117 390 133 547
rect 145 390 161 602
rect 172 390 188 602
rect 199 390 219 602
rect 230 390 246 680
rect 257 390 273 680
rect 284 390 300 680
rect 311 390 327 680
<< psubstratetap >>
rect 9 70 25 86
rect 37 70 53 86
rect 65 70 81 86
rect 93 70 109 86
rect 121 70 137 86
rect 149 70 165 86
rect 177 70 193 86
rect 205 70 221 86
rect 233 70 250 86
rect 262 70 278 86
rect 290 70 306 86
rect 318 70 334 86
<< nsubstratetap >>
rect 9 712 25 728
rect 37 712 53 728
rect 65 712 81 728
rect 93 712 109 728
rect 121 712 137 728
rect 149 712 165 728
rect 177 712 193 728
rect 205 712 221 728
rect 233 712 250 728
rect 262 712 278 728
rect 290 712 306 728
rect 318 712 334 728
<< metal1 >>
rect 3 766 340 776
rect 3 742 340 752
rect 3 712 9 728
rect 25 712 37 728
rect 53 712 65 728
rect 81 712 93 728
rect 109 712 121 728
rect 137 712 149 728
rect 165 712 177 728
rect 193 712 205 728
rect 221 712 233 728
rect 250 712 262 728
rect 278 712 290 728
rect 306 712 318 728
rect 334 712 340 728
rect 3 703 340 712
rect 35 448 51 703
rect 90 547 106 703
rect 145 602 161 703
rect 199 680 219 703
rect 257 680 273 703
rect 311 680 327 703
rect 199 602 202 680
rect 3 363 42 373
rect 68 373 78 390
rect 68 363 97 373
rect 68 350 78 363
rect 123 374 133 390
rect 123 364 152 374
rect 123 350 133 364
rect 178 374 188 390
rect 178 364 210 374
rect 178 350 188 364
rect 236 375 246 390
rect 290 375 300 390
rect 236 365 340 375
rect 236 350 246 365
rect 35 95 51 330
rect 90 95 106 296
rect 145 95 161 204
rect 203 95 219 150
rect 257 95 273 150
rect 3 86 340 95
rect 3 70 9 86
rect 25 70 37 86
rect 53 70 65 86
rect 81 70 93 86
rect 109 70 121 86
rect 137 70 149 86
rect 165 70 177 86
rect 193 70 205 86
rect 221 70 233 86
rect 250 70 262 86
rect 278 70 290 86
rect 306 70 318 86
rect 334 70 340 86
rect 3 47 340 57
rect 3 24 340 34
rect 3 1 340 11
<< end >>
