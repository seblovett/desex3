magic
tech c035u
timestamp 1385033586
<< nwell >>
rect 230 532 1527 744
rect 230 497 1415 532
rect 230 496 1399 497
rect 352 404 669 496
rect 717 404 1034 496
rect 1082 404 1399 496
rect 405 403 451 404
rect 770 403 816 404
rect 1135 403 1181 404
<< polysilicon >>
rect 563 694 570 702
rect 590 694 597 702
rect 617 694 624 702
rect 644 694 651 702
rect 928 694 935 702
rect 955 694 962 702
rect 982 694 989 702
rect 1009 694 1016 702
rect 1293 694 1300 702
rect 1320 694 1327 702
rect 1347 694 1354 702
rect 1374 694 1381 702
rect 480 616 487 624
rect 507 616 514 624
rect 425 561 432 569
rect 370 462 377 470
rect 845 616 852 624
rect 872 616 879 624
rect 790 561 797 569
rect 735 462 742 470
rect 1210 616 1217 624
rect 1237 616 1244 624
rect 1155 561 1162 569
rect 1100 462 1107 470
rect 1479 645 1481 661
rect 1474 600 1481 645
rect 1474 504 1481 552
rect 1474 466 1481 474
rect 370 390 377 404
rect 425 390 432 404
rect 480 391 487 404
rect 375 374 377 390
rect 430 374 432 390
rect 485 387 487 391
rect 507 387 514 404
rect 563 391 570 404
rect 485 380 514 387
rect 485 375 487 380
rect 568 387 570 391
rect 590 387 597 404
rect 617 387 624 404
rect 644 387 651 404
rect 735 390 742 404
rect 790 390 797 404
rect 845 391 852 404
rect 568 380 651 387
rect 568 375 570 380
rect 370 364 377 374
rect 425 364 432 374
rect 480 364 487 375
rect 563 364 570 375
rect 590 364 597 380
rect 740 374 742 390
rect 795 374 797 390
rect 850 387 852 391
rect 872 387 879 404
rect 928 391 935 404
rect 850 380 879 387
rect 850 375 852 380
rect 933 387 935 391
rect 955 387 962 404
rect 982 387 989 404
rect 1009 387 1016 404
rect 1100 390 1107 404
rect 1155 390 1162 404
rect 1210 391 1217 404
rect 933 380 1016 387
rect 933 375 935 380
rect 735 364 742 374
rect 790 364 797 374
rect 845 364 852 375
rect 928 364 935 375
rect 955 364 962 380
rect 1105 374 1107 390
rect 1160 374 1162 390
rect 1215 387 1217 391
rect 1237 387 1244 404
rect 1293 391 1300 404
rect 1215 380 1244 387
rect 1215 375 1217 380
rect 1298 387 1300 391
rect 1320 387 1327 404
rect 1347 387 1354 404
rect 1374 387 1381 404
rect 1298 380 1381 387
rect 1298 375 1300 380
rect 1100 364 1107 374
rect 1155 364 1162 374
rect 1210 364 1217 375
rect 1293 364 1300 375
rect 1320 364 1327 380
rect 370 336 377 344
rect 425 302 432 310
rect 480 210 487 218
rect 735 336 742 344
rect 790 302 797 310
rect 845 210 852 218
rect 1100 336 1107 344
rect 1155 302 1162 310
rect 1210 210 1217 218
rect 563 156 570 164
rect 590 156 597 164
rect 928 156 935 164
rect 955 156 962 164
rect 1293 156 1300 164
rect 1320 156 1327 164
<< ndiffusion >>
rect 1472 474 1474 504
rect 1481 474 1483 504
rect 368 344 370 364
rect 377 344 379 364
rect 423 310 425 364
rect 432 310 434 364
rect 478 218 480 364
rect 487 218 489 364
rect 561 164 563 364
rect 570 164 572 364
rect 588 164 590 364
rect 597 164 599 364
rect 733 344 735 364
rect 742 344 744 364
rect 788 310 790 364
rect 797 310 799 364
rect 843 218 845 364
rect 852 218 854 364
rect 926 164 928 364
rect 935 164 937 364
rect 953 164 955 364
rect 962 164 964 364
rect 1098 344 1100 364
rect 1107 344 1109 364
rect 1153 310 1155 364
rect 1162 310 1164 364
rect 1208 218 1210 364
rect 1217 218 1219 364
rect 1291 164 1293 364
rect 1300 164 1302 364
rect 1318 164 1320 364
rect 1327 164 1329 364
<< pdiffusion >>
rect 368 404 370 462
rect 377 404 379 462
rect 423 404 425 561
rect 432 404 434 561
rect 478 404 480 616
rect 487 404 489 616
rect 505 404 507 616
rect 514 404 516 616
rect 561 404 563 694
rect 570 404 572 694
rect 588 404 590 694
rect 597 404 599 694
rect 615 404 617 694
rect 624 404 626 694
rect 642 404 644 694
rect 651 404 653 694
rect 733 404 735 462
rect 742 404 744 462
rect 788 404 790 561
rect 797 404 799 561
rect 843 404 845 616
rect 852 404 854 616
rect 870 404 872 616
rect 879 404 881 616
rect 926 404 928 694
rect 935 404 937 694
rect 953 404 955 694
rect 962 404 964 694
rect 980 404 982 694
rect 989 404 991 694
rect 1007 404 1009 694
rect 1016 404 1018 694
rect 1098 404 1100 462
rect 1107 404 1109 462
rect 1153 404 1155 561
rect 1162 404 1164 561
rect 1208 404 1210 616
rect 1217 404 1219 616
rect 1235 404 1237 616
rect 1244 404 1246 616
rect 1291 404 1293 694
rect 1300 404 1302 694
rect 1318 404 1320 694
rect 1327 404 1329 694
rect 1345 404 1347 694
rect 1354 404 1356 694
rect 1372 404 1374 694
rect 1381 404 1383 694
rect 1472 552 1474 600
rect 1481 552 1483 600
<< pohmic >>
rect 352 84 354 94
rect 370 84 382 94
rect 398 84 410 94
rect 426 84 438 94
rect 454 84 466 94
rect 482 84 494 94
rect 510 84 522 94
rect 538 84 550 94
rect 567 84 579 94
rect 595 84 607 94
rect 623 84 635 94
rect 651 84 663 94
rect 679 84 691 94
rect 707 84 719 94
rect 735 84 747 94
rect 763 84 775 94
rect 791 84 803 94
rect 819 84 831 94
rect 847 84 859 94
rect 875 84 887 94
rect 903 84 915 94
rect 932 84 944 94
rect 960 84 972 94
rect 988 84 1000 94
rect 1016 84 1028 94
rect 1044 84 1056 94
rect 1072 84 1084 94
rect 1100 84 1112 94
rect 1128 84 1140 94
rect 1156 84 1168 94
rect 1184 84 1196 94
rect 1212 84 1224 94
rect 1240 84 1252 94
rect 1268 84 1280 94
rect 1297 84 1309 94
rect 1325 84 1337 94
rect 1353 84 1365 94
rect 1381 84 1393 94
rect 1409 84 1421 94
rect 1437 84 1449 94
rect 1465 84 1477 94
rect 1493 84 1505 94
rect 1521 84 1527 94
<< nohmic >>
rect 230 734 242 744
rect 258 734 270 744
rect 286 734 298 744
rect 314 734 326 744
rect 342 734 354 744
rect 370 734 382 744
rect 398 734 410 744
rect 426 734 438 744
rect 454 734 466 744
rect 482 734 494 744
rect 510 734 522 744
rect 538 734 550 744
rect 567 734 579 744
rect 595 734 607 744
rect 623 734 635 744
rect 651 734 663 744
rect 679 734 691 744
rect 707 734 719 744
rect 735 734 747 744
rect 763 734 775 744
rect 791 734 803 744
rect 819 734 831 744
rect 847 734 859 744
rect 875 734 887 744
rect 903 734 915 744
rect 932 734 944 744
rect 960 734 972 744
rect 988 734 1000 744
rect 1016 734 1028 744
rect 1044 734 1056 744
rect 1072 734 1084 744
rect 1100 734 1112 744
rect 1128 734 1140 744
rect 1156 734 1168 744
rect 1184 734 1196 744
rect 1212 734 1224 744
rect 1240 734 1252 744
rect 1268 734 1280 744
rect 1297 734 1309 744
rect 1325 734 1337 744
rect 1353 734 1365 744
rect 1381 734 1393 744
rect 1409 734 1421 744
rect 1437 734 1449 744
rect 1465 734 1477 744
rect 1493 734 1505 744
rect 1521 734 1527 744
<< ntransistor >>
rect 1474 474 1481 504
rect 370 344 377 364
rect 425 310 432 364
rect 480 218 487 364
rect 563 164 570 364
rect 590 164 597 364
rect 735 344 742 364
rect 790 310 797 364
rect 845 218 852 364
rect 928 164 935 364
rect 955 164 962 364
rect 1100 344 1107 364
rect 1155 310 1162 364
rect 1210 218 1217 364
rect 1293 164 1300 364
rect 1320 164 1327 364
<< ptransistor >>
rect 370 404 377 462
rect 425 404 432 561
rect 480 404 487 616
rect 507 404 514 616
rect 563 404 570 694
rect 590 404 597 694
rect 617 404 624 694
rect 644 404 651 694
rect 735 404 742 462
rect 790 404 797 561
rect 845 404 852 616
rect 872 404 879 616
rect 928 404 935 694
rect 955 404 962 694
rect 982 404 989 694
rect 1009 404 1016 694
rect 1100 404 1107 462
rect 1155 404 1162 561
rect 1210 404 1217 616
rect 1237 404 1244 616
rect 1293 404 1300 694
rect 1320 404 1327 694
rect 1347 404 1354 694
rect 1374 404 1381 694
rect 1474 552 1481 600
<< polycontact >>
rect 1463 645 1479 661
rect 359 374 375 390
rect 414 374 430 390
rect 469 375 485 391
rect 552 375 568 391
rect 724 374 740 390
rect 779 374 795 390
rect 834 375 850 391
rect 917 375 933 391
rect 1089 374 1105 390
rect 1144 374 1160 390
rect 1199 375 1215 391
rect 1282 375 1298 391
<< ndiffcontact >>
rect 1456 474 1472 504
rect 1483 474 1499 504
rect 352 344 368 364
rect 379 344 395 364
rect 407 310 423 364
rect 434 310 450 364
rect 462 218 478 364
rect 489 218 505 364
rect 545 164 561 364
rect 572 164 588 364
rect 599 164 615 364
rect 717 344 733 364
rect 744 344 760 364
rect 772 310 788 364
rect 799 310 815 364
rect 827 218 843 364
rect 854 218 870 364
rect 910 164 926 364
rect 937 164 953 364
rect 964 164 980 364
rect 1082 344 1098 364
rect 1109 344 1125 364
rect 1137 310 1153 364
rect 1164 310 1180 364
rect 1192 218 1208 364
rect 1219 218 1235 364
rect 1275 164 1291 364
rect 1302 164 1318 364
rect 1329 164 1345 364
<< pdiffcontact >>
rect 352 404 368 462
rect 379 404 395 462
rect 407 404 423 561
rect 434 404 450 561
rect 462 404 478 616
rect 489 404 505 616
rect 516 404 532 616
rect 545 404 561 694
rect 572 404 588 694
rect 599 404 615 694
rect 626 404 642 694
rect 653 404 669 694
rect 717 404 733 462
rect 744 404 760 462
rect 772 404 788 561
rect 799 404 815 561
rect 827 404 843 616
rect 854 404 870 616
rect 881 404 897 616
rect 910 404 926 694
rect 937 404 953 694
rect 964 404 980 694
rect 991 404 1007 694
rect 1018 404 1034 694
rect 1082 404 1098 462
rect 1109 404 1125 462
rect 1137 404 1153 561
rect 1164 404 1180 561
rect 1192 404 1208 616
rect 1219 404 1235 616
rect 1246 404 1262 616
rect 1275 404 1291 694
rect 1302 404 1318 694
rect 1329 404 1345 694
rect 1356 404 1372 694
rect 1383 404 1399 694
rect 1456 552 1472 600
rect 1483 552 1499 600
<< psubstratetap >>
rect 354 84 370 100
rect 382 84 398 100
rect 410 84 426 100
rect 438 84 454 100
rect 466 84 482 100
rect 494 84 510 100
rect 522 84 538 100
rect 550 84 567 100
rect 579 84 595 100
rect 607 84 623 100
rect 635 84 651 100
rect 663 84 679 100
rect 691 84 707 100
rect 719 84 735 100
rect 747 84 763 100
rect 775 84 791 100
rect 803 84 819 100
rect 831 84 847 100
rect 859 84 875 100
rect 887 84 903 100
rect 915 84 932 100
rect 944 84 960 100
rect 972 84 988 100
rect 1000 84 1016 100
rect 1028 84 1044 100
rect 1056 84 1072 100
rect 1084 84 1100 100
rect 1112 84 1128 100
rect 1140 84 1156 100
rect 1168 84 1184 100
rect 1196 84 1212 100
rect 1224 84 1240 100
rect 1252 84 1268 100
rect 1280 84 1297 100
rect 1309 84 1325 100
rect 1337 84 1353 100
rect 1365 84 1381 100
rect 1393 84 1409 100
rect 1421 84 1437 100
rect 1449 84 1465 100
rect 1477 84 1493 100
rect 1505 84 1521 100
<< nsubstratetap >>
rect 242 728 258 744
rect 270 728 286 744
rect 298 728 314 744
rect 326 728 342 744
rect 354 728 370 744
rect 382 728 398 744
rect 410 728 426 744
rect 438 728 454 744
rect 466 728 482 744
rect 494 728 510 744
rect 522 728 538 744
rect 550 728 567 744
rect 579 728 595 744
rect 607 728 623 744
rect 635 728 651 744
rect 663 728 679 744
rect 691 728 707 744
rect 719 728 735 744
rect 747 728 763 744
rect 775 728 791 744
rect 803 728 819 744
rect 831 728 847 744
rect 859 728 875 744
rect 887 728 903 744
rect 915 728 932 744
rect 944 728 960 744
rect 972 728 988 744
rect 1000 728 1016 744
rect 1028 728 1044 744
rect 1056 728 1072 744
rect 1084 728 1100 744
rect 1112 728 1128 744
rect 1140 728 1156 744
rect 1168 728 1184 744
rect 1196 728 1212 744
rect 1224 728 1240 744
rect 1252 728 1268 744
rect 1280 728 1297 744
rect 1309 728 1325 744
rect 1337 728 1353 744
rect 1365 728 1381 744
rect 1393 728 1409 744
rect 1421 728 1437 744
rect 1449 728 1465 744
rect 1477 728 1493 744
rect 1505 728 1521 744
<< metal1 >>
rect 264 780 1441 790
rect 1485 780 1527 790
rect 264 757 1527 767
rect 228 728 242 744
rect 258 728 270 744
rect 286 728 298 744
rect 314 728 326 744
rect 342 728 354 744
rect 370 728 382 744
rect 398 728 410 744
rect 426 728 438 744
rect 454 728 466 744
rect 482 728 494 744
rect 510 728 522 744
rect 538 728 550 744
rect 567 728 579 744
rect 595 728 607 744
rect 623 728 635 744
rect 651 728 663 744
rect 679 728 691 744
rect 707 728 719 744
rect 735 728 747 744
rect 763 728 775 744
rect 791 728 803 744
rect 819 728 831 744
rect 847 728 859 744
rect 875 728 887 744
rect 903 728 915 744
rect 932 728 944 744
rect 960 728 972 744
rect 988 728 1000 744
rect 1016 728 1028 744
rect 1044 728 1056 744
rect 1072 728 1084 744
rect 1100 728 1112 744
rect 1128 728 1140 744
rect 1156 728 1168 744
rect 1184 728 1196 744
rect 1212 728 1224 744
rect 1240 728 1252 744
rect 1268 728 1280 744
rect 1297 728 1309 744
rect 1325 728 1337 744
rect 1353 728 1365 744
rect 1381 728 1393 744
rect 1409 728 1421 744
rect 1437 728 1449 744
rect 1465 728 1477 744
rect 1493 728 1505 744
rect 1521 728 1527 744
rect 228 719 1527 728
rect 352 462 368 719
rect 407 561 423 719
rect 462 616 478 719
rect 516 616 532 719
rect 545 694 561 719
rect 599 694 615 719
rect 653 694 669 719
rect 717 462 733 719
rect 772 561 788 719
rect 827 616 843 719
rect 881 616 897 719
rect 910 694 926 719
rect 964 694 980 719
rect 1018 694 1034 719
rect 1082 462 1098 719
rect 1137 561 1153 719
rect 1192 616 1208 719
rect 1246 616 1262 719
rect 1275 694 1291 719
rect 1329 694 1345 719
rect 1383 694 1399 719
rect 1465 661 1479 667
rect 1489 600 1499 719
rect 1456 504 1466 552
rect 312 377 359 387
rect 385 387 395 404
rect 385 377 414 387
rect 385 364 395 377
rect 440 388 450 404
rect 440 378 469 388
rect 440 364 450 378
rect 495 388 505 404
rect 495 378 552 388
rect 495 364 505 378
rect 578 389 588 404
rect 632 391 642 404
rect 578 379 630 389
rect 578 364 588 379
rect 713 377 724 387
rect 750 387 760 404
rect 750 377 779 387
rect 750 364 760 377
rect 805 388 815 404
rect 805 378 834 388
rect 805 364 815 378
rect 860 388 870 404
rect 860 378 917 388
rect 860 364 870 378
rect 943 389 953 404
rect 997 391 1007 404
rect 943 379 993 389
rect 943 364 953 379
rect 1079 377 1089 387
rect 1115 387 1125 404
rect 1115 377 1144 387
rect 1115 364 1125 377
rect 1170 388 1180 404
rect 1170 378 1199 388
rect 1170 364 1180 378
rect 1225 388 1235 404
rect 1225 378 1282 388
rect 1225 364 1235 378
rect 1308 389 1318 404
rect 1362 391 1372 404
rect 1308 379 1356 389
rect 1308 364 1318 379
rect 1370 389 1372 391
rect 1370 379 1415 389
rect 352 109 368 344
rect 407 109 423 310
rect 462 109 478 218
rect 545 109 561 164
rect 599 109 615 164
rect 717 109 733 344
rect 772 109 788 310
rect 827 109 843 218
rect 910 109 926 164
rect 964 109 980 164
rect 1082 109 1098 344
rect 1137 109 1153 310
rect 1192 109 1208 218
rect 1275 109 1291 164
rect 1329 109 1345 164
rect 1483 109 1493 474
rect 352 100 1527 109
rect 352 84 354 100
rect 370 84 382 100
rect 398 84 410 100
rect 426 84 438 100
rect 454 84 466 100
rect 482 84 494 100
rect 510 84 522 100
rect 538 84 550 100
rect 567 84 579 100
rect 595 84 607 100
rect 623 84 635 100
rect 651 84 663 100
rect 679 84 691 100
rect 707 84 719 100
rect 735 84 747 100
rect 763 84 775 100
rect 791 84 803 100
rect 819 84 831 100
rect 847 84 859 100
rect 875 84 887 100
rect 903 84 915 100
rect 932 84 944 100
rect 960 84 972 100
rect 988 84 1000 100
rect 1016 84 1028 100
rect 1044 84 1056 100
rect 1072 84 1084 100
rect 1100 84 1112 100
rect 1128 84 1140 100
rect 1156 84 1168 100
rect 1184 84 1196 100
rect 1212 84 1224 100
rect 1240 84 1252 100
rect 1268 84 1280 100
rect 1297 84 1309 100
rect 1325 84 1337 100
rect 1353 84 1365 100
rect 1381 84 1393 100
rect 1409 84 1421 100
rect 1437 84 1449 100
rect 1465 84 1477 100
rect 1493 84 1505 100
rect 1521 84 1527 100
rect 645 61 1527 71
rect 288 38 699 48
rect 1008 38 1527 48
rect 336 15 1064 25
rect 1371 15 1527 25
<< m2contact >>
rect 250 779 264 793
rect 1441 779 1455 793
rect 1471 779 1485 793
rect 250 755 264 769
rect 28 719 228 744
rect 1465 667 1479 681
rect 1442 586 1456 600
rect 298 375 312 389
rect 630 377 644 391
rect 699 375 713 389
rect 993 377 1007 391
rect 1065 375 1079 389
rect 1356 377 1370 391
rect 631 59 645 73
rect 274 37 288 51
rect 699 36 713 50
rect 994 36 1008 50
rect 322 13 336 27
rect 1064 13 1078 27
rect 1357 13 1371 27
<< metal2 >>
rect 28 744 228 798
rect 251 793 263 798
rect 28 8 228 719
rect 251 8 263 755
rect 275 51 287 798
rect 299 389 311 798
rect 275 8 287 37
rect 299 8 311 375
rect 323 27 335 798
rect 1443 600 1455 779
rect 1471 681 1483 779
rect 1479 667 1483 681
rect 632 73 644 377
rect 700 50 712 375
rect 995 50 1007 377
rect 1065 27 1077 375
rect 1358 27 1370 377
rect 323 8 335 13
<< labels >>
rlabel metal1 1527 780 1527 790 7 nSDO
rlabel metal1 1527 757 1527 767 7 SDI
rlabel metal1 1527 719 1527 744 7 Vdd!
rlabel metal1 1527 84 1527 109 7 GND!
rlabel metal1 1527 61 1527 71 7 ClockOut
rlabel metal1 1527 38 1527 48 7 TestOut
rlabel metal1 1527 15 1527 25 7 nResetOut
rlabel metal2 275 8 287 8 1 Test
rlabel metal2 299 8 311 8 1 Clock
rlabel metal2 28 8 228 8 1 Vdd!
rlabel metal2 323 8 335 8 1 nReset
rlabel metal2 251 8 263 8 1 SDI
rlabel metal2 323 798 335 798 5 nReset
rlabel metal2 299 798 311 798 5 Clock
rlabel metal2 275 798 287 798 5 Test
rlabel metal2 251 798 263 798 5 SDO
rlabel metal2 28 798 228 798 5 Vdd!
<< end >>
