magic
tech c035u
timestamp 1384526628
<< nwell >>
rect 324 207 1929 419
<< polysilicon >>
rect 433 384 440 392
rect 928 384 935 392
rect 1417 384 1424 392
rect 378 285 385 293
rect 488 368 495 376
rect 515 368 522 376
rect 542 368 549 376
rect 597 372 604 380
rect 624 372 631 380
rect 651 372 658 380
rect 678 372 685 380
rect 705 372 712 380
rect 732 372 739 380
rect 759 372 766 380
rect 786 372 793 380
rect 873 285 880 293
rect 983 368 990 376
rect 1010 368 1017 376
rect 1037 368 1044 376
rect 1092 372 1099 380
rect 1119 372 1126 380
rect 1146 372 1153 380
rect 1173 372 1180 380
rect 1200 372 1207 380
rect 1227 372 1234 380
rect 1254 372 1261 380
rect 1281 372 1288 380
rect 1362 285 1369 293
rect 1472 368 1479 376
rect 1499 368 1506 376
rect 1526 368 1533 376
rect 1581 372 1588 380
rect 1608 372 1615 380
rect 1635 372 1642 380
rect 1662 372 1669 380
rect 1689 372 1696 380
rect 1716 372 1723 380
rect 1743 372 1750 380
rect 1770 372 1777 380
rect 1869 348 1871 364
rect 1864 275 1871 348
rect 378 213 385 227
rect 433 213 440 227
rect 488 213 495 227
rect 383 197 385 213
rect 438 197 440 213
rect 493 208 495 213
rect 515 208 522 227
rect 542 208 549 227
rect 597 213 604 227
rect 493 201 549 208
rect 493 197 495 201
rect 378 187 385 197
rect 433 187 440 197
rect 488 187 495 197
rect 515 187 522 201
rect 602 208 604 213
rect 624 208 631 227
rect 651 208 658 227
rect 678 208 685 227
rect 705 208 712 227
rect 732 208 739 227
rect 759 208 766 227
rect 786 210 793 227
rect 873 213 880 227
rect 928 213 935 227
rect 983 213 990 227
rect 784 208 793 210
rect 602 201 793 208
rect 602 197 604 201
rect 597 187 604 197
rect 624 187 631 201
rect 651 187 658 201
rect 678 187 685 201
rect 705 187 712 201
rect 732 187 739 201
rect 759 187 766 201
rect 786 187 793 201
rect 878 197 880 213
rect 933 197 935 213
rect 988 208 990 213
rect 1010 208 1017 227
rect 1037 208 1044 227
rect 1092 213 1099 227
rect 988 201 1044 208
rect 988 197 990 201
rect 873 187 880 197
rect 928 187 935 197
rect 983 187 990 197
rect 1010 187 1017 201
rect 1097 208 1099 213
rect 1119 208 1126 227
rect 1146 208 1153 227
rect 1173 208 1180 227
rect 1200 208 1207 227
rect 1227 208 1234 227
rect 1254 208 1261 227
rect 1281 210 1288 227
rect 1362 213 1369 227
rect 1417 213 1424 227
rect 1472 213 1479 227
rect 1279 208 1288 210
rect 1097 201 1288 208
rect 1097 197 1099 201
rect 1092 187 1099 197
rect 1119 187 1126 201
rect 1146 187 1153 201
rect 1173 187 1180 201
rect 1200 187 1207 201
rect 1227 187 1234 201
rect 1254 187 1261 201
rect 1281 187 1288 201
rect 1367 197 1369 213
rect 1422 197 1424 213
rect 1477 208 1479 213
rect 1499 208 1506 227
rect 1526 208 1533 227
rect 1581 213 1588 227
rect 1477 201 1533 208
rect 1477 197 1479 201
rect 1362 187 1369 197
rect 1417 187 1424 197
rect 1472 187 1479 197
rect 1499 187 1506 201
rect 1586 208 1588 213
rect 1608 208 1615 227
rect 1635 208 1642 227
rect 1662 208 1669 227
rect 1689 208 1696 227
rect 1716 208 1723 227
rect 1743 208 1750 227
rect 1770 210 1777 227
rect 1768 208 1777 210
rect 1586 201 1777 208
rect 1586 197 1588 201
rect 1581 187 1588 197
rect 1608 187 1615 201
rect 1635 187 1642 201
rect 1662 187 1669 201
rect 1689 187 1696 201
rect 1716 187 1723 201
rect 1743 187 1750 201
rect 1770 187 1777 201
rect 1864 187 1871 227
rect 378 159 385 167
rect 433 125 440 133
rect 873 159 880 167
rect 597 129 604 137
rect 624 129 631 137
rect 651 129 658 137
rect 678 129 685 137
rect 705 129 712 137
rect 732 129 739 137
rect 759 129 766 137
rect 786 129 793 137
rect 928 125 935 133
rect 1362 159 1369 167
rect 1092 129 1099 137
rect 1119 129 1126 137
rect 1146 129 1153 137
rect 1173 129 1180 137
rect 1200 129 1207 137
rect 1227 129 1234 137
rect 1254 129 1261 137
rect 1281 129 1288 137
rect 1417 125 1424 133
rect 1864 149 1871 157
rect 1581 129 1588 137
rect 1608 129 1615 137
rect 1635 129 1642 137
rect 1662 129 1669 137
rect 1689 129 1696 137
rect 1716 129 1723 137
rect 1743 129 1750 137
rect 1770 129 1777 137
rect 488 106 495 114
rect 515 106 522 114
rect 983 106 990 114
rect 1010 106 1017 114
rect 1472 106 1479 114
rect 1499 106 1506 114
<< ndiffusion >>
rect 376 167 378 187
rect 385 167 387 187
rect 431 133 433 187
rect 440 133 442 187
rect 486 114 488 187
rect 495 114 497 187
rect 513 114 515 187
rect 522 114 524 187
rect 595 137 597 187
rect 604 137 606 187
rect 622 137 624 187
rect 631 137 633 187
rect 649 137 651 187
rect 658 137 660 187
rect 676 137 678 187
rect 685 137 687 187
rect 703 137 705 187
rect 712 137 714 187
rect 730 137 732 187
rect 739 137 741 187
rect 757 137 759 187
rect 766 137 768 187
rect 784 137 786 187
rect 793 137 795 187
rect 871 167 873 187
rect 880 167 882 187
rect 926 133 928 187
rect 935 133 937 187
rect 981 114 983 187
rect 990 114 992 187
rect 1008 114 1010 187
rect 1017 114 1019 187
rect 1090 137 1092 187
rect 1099 137 1101 187
rect 1117 137 1119 187
rect 1126 137 1128 187
rect 1144 137 1146 187
rect 1153 137 1155 187
rect 1171 137 1173 187
rect 1180 137 1182 187
rect 1198 137 1200 187
rect 1207 137 1209 187
rect 1225 137 1227 187
rect 1234 137 1236 187
rect 1252 137 1254 187
rect 1261 137 1263 187
rect 1279 137 1281 187
rect 1288 137 1290 187
rect 1360 167 1362 187
rect 1369 167 1371 187
rect 1415 133 1417 187
rect 1424 133 1426 187
rect 1470 114 1472 187
rect 1479 114 1481 187
rect 1497 114 1499 187
rect 1506 114 1508 187
rect 1579 137 1581 187
rect 1588 137 1590 187
rect 1606 137 1608 187
rect 1615 137 1617 187
rect 1633 137 1635 187
rect 1642 137 1644 187
rect 1660 137 1662 187
rect 1669 137 1671 187
rect 1687 137 1689 187
rect 1696 137 1698 187
rect 1714 137 1716 187
rect 1723 137 1725 187
rect 1741 137 1743 187
rect 1750 137 1752 187
rect 1768 137 1770 187
rect 1777 137 1779 187
rect 1862 157 1864 187
rect 1871 157 1873 187
<< pdiffusion >>
rect 376 227 378 285
rect 385 227 387 285
rect 431 227 433 384
rect 440 227 442 384
rect 486 227 488 368
rect 495 227 497 368
rect 513 227 515 368
rect 522 227 524 368
rect 540 227 542 368
rect 549 227 551 368
rect 595 227 597 372
rect 604 227 606 372
rect 622 227 624 372
rect 631 227 633 372
rect 649 227 651 372
rect 658 227 660 372
rect 676 227 678 372
rect 685 227 687 372
rect 703 227 705 372
rect 712 227 714 372
rect 730 227 732 372
rect 739 227 741 372
rect 757 227 759 372
rect 766 227 768 372
rect 784 227 786 372
rect 793 227 795 372
rect 871 227 873 285
rect 880 227 882 285
rect 926 227 928 384
rect 935 227 937 384
rect 981 227 983 368
rect 990 227 992 368
rect 1008 227 1010 368
rect 1017 227 1019 368
rect 1035 227 1037 368
rect 1044 227 1046 368
rect 1090 227 1092 372
rect 1099 227 1101 372
rect 1117 227 1119 372
rect 1126 227 1128 372
rect 1144 227 1146 372
rect 1153 227 1155 372
rect 1171 227 1173 372
rect 1180 227 1182 372
rect 1198 227 1200 372
rect 1207 227 1209 372
rect 1225 227 1227 372
rect 1234 227 1236 372
rect 1252 227 1254 372
rect 1261 227 1263 372
rect 1279 227 1281 372
rect 1288 227 1290 372
rect 1360 227 1362 285
rect 1369 227 1371 285
rect 1415 227 1417 384
rect 1424 227 1426 384
rect 1470 227 1472 368
rect 1479 227 1481 368
rect 1497 227 1499 368
rect 1506 227 1508 368
rect 1524 227 1526 368
rect 1533 227 1535 368
rect 1579 227 1581 372
rect 1588 227 1590 372
rect 1606 227 1608 372
rect 1615 227 1617 372
rect 1633 227 1635 372
rect 1642 227 1644 372
rect 1660 227 1662 372
rect 1669 227 1671 372
rect 1687 227 1689 372
rect 1696 227 1698 372
rect 1714 227 1716 372
rect 1723 227 1725 372
rect 1741 227 1743 372
rect 1750 227 1752 372
rect 1768 227 1770 372
rect 1777 227 1779 372
rect 1862 227 1864 275
rect 1871 227 1873 275
<< nohmic >>
rect 324 409 1929 419
<< ntransistor >>
rect 378 167 385 187
rect 433 133 440 187
rect 488 114 495 187
rect 515 114 522 187
rect 597 137 604 187
rect 624 137 631 187
rect 651 137 658 187
rect 678 137 685 187
rect 705 137 712 187
rect 732 137 739 187
rect 759 137 766 187
rect 786 137 793 187
rect 873 167 880 187
rect 928 133 935 187
rect 983 114 990 187
rect 1010 114 1017 187
rect 1092 137 1099 187
rect 1119 137 1126 187
rect 1146 137 1153 187
rect 1173 137 1180 187
rect 1200 137 1207 187
rect 1227 137 1234 187
rect 1254 137 1261 187
rect 1281 137 1288 187
rect 1362 167 1369 187
rect 1417 133 1424 187
rect 1472 114 1479 187
rect 1499 114 1506 187
rect 1581 137 1588 187
rect 1608 137 1615 187
rect 1635 137 1642 187
rect 1662 137 1669 187
rect 1689 137 1696 187
rect 1716 137 1723 187
rect 1743 137 1750 187
rect 1770 137 1777 187
rect 1864 157 1871 187
<< ptransistor >>
rect 378 227 385 285
rect 433 227 440 384
rect 488 227 495 368
rect 515 227 522 368
rect 542 227 549 368
rect 597 227 604 372
rect 624 227 631 372
rect 651 227 658 372
rect 678 227 685 372
rect 705 227 712 372
rect 732 227 739 372
rect 759 227 766 372
rect 786 227 793 372
rect 873 227 880 285
rect 928 227 935 384
rect 983 227 990 368
rect 1010 227 1017 368
rect 1037 227 1044 368
rect 1092 227 1099 372
rect 1119 227 1126 372
rect 1146 227 1153 372
rect 1173 227 1180 372
rect 1200 227 1207 372
rect 1227 227 1234 372
rect 1254 227 1261 372
rect 1281 227 1288 372
rect 1362 227 1369 285
rect 1417 227 1424 384
rect 1472 227 1479 368
rect 1499 227 1506 368
rect 1526 227 1533 368
rect 1581 227 1588 372
rect 1608 227 1615 372
rect 1635 227 1642 372
rect 1662 227 1669 372
rect 1689 227 1696 372
rect 1716 227 1723 372
rect 1743 227 1750 372
rect 1770 227 1777 372
rect 1864 227 1871 275
<< polycontact >>
rect 1853 348 1869 364
rect 367 197 383 213
rect 422 197 438 213
rect 477 197 493 213
rect 586 197 602 213
rect 862 197 878 213
rect 917 197 933 213
rect 972 197 988 213
rect 1081 197 1097 213
rect 1351 197 1367 213
rect 1406 197 1422 213
rect 1461 197 1477 213
rect 1570 197 1586 213
<< ndiffcontact >>
rect 360 167 376 187
rect 387 167 403 187
rect 415 133 431 187
rect 442 133 458 187
rect 470 114 486 187
rect 497 114 513 187
rect 524 114 540 187
rect 579 137 595 187
rect 606 137 622 187
rect 633 137 649 187
rect 660 137 676 187
rect 687 137 703 187
rect 714 137 730 187
rect 741 137 757 187
rect 768 137 784 187
rect 795 137 811 187
rect 855 167 871 187
rect 882 167 898 187
rect 910 133 926 187
rect 937 133 953 187
rect 965 114 981 187
rect 992 114 1008 187
rect 1019 114 1035 187
rect 1074 137 1090 187
rect 1101 137 1117 187
rect 1128 137 1144 187
rect 1155 137 1171 187
rect 1182 137 1198 187
rect 1209 137 1225 187
rect 1236 137 1252 187
rect 1263 137 1279 187
rect 1290 137 1306 187
rect 1344 167 1360 187
rect 1371 167 1387 187
rect 1399 133 1415 187
rect 1426 133 1442 187
rect 1454 114 1470 187
rect 1481 114 1497 187
rect 1508 114 1524 187
rect 1563 137 1579 187
rect 1590 137 1606 187
rect 1617 137 1633 187
rect 1644 137 1660 187
rect 1671 137 1687 187
rect 1698 137 1714 187
rect 1725 137 1741 187
rect 1752 137 1768 187
rect 1779 137 1795 187
rect 1846 157 1862 187
rect 1873 157 1889 187
<< pdiffcontact >>
rect 360 227 376 285
rect 387 227 403 285
rect 415 227 431 384
rect 442 227 458 384
rect 470 227 486 368
rect 497 227 513 368
rect 524 227 540 368
rect 551 227 567 368
rect 579 227 595 372
rect 606 227 622 372
rect 633 227 649 372
rect 660 227 676 372
rect 687 227 703 372
rect 714 227 730 372
rect 741 227 757 372
rect 768 227 784 372
rect 795 227 811 372
rect 855 227 871 285
rect 882 227 898 285
rect 910 227 926 384
rect 937 227 953 384
rect 965 227 981 368
rect 992 227 1008 368
rect 1019 227 1035 368
rect 1046 227 1062 368
rect 1074 227 1090 372
rect 1101 227 1117 372
rect 1128 227 1144 372
rect 1155 227 1171 372
rect 1182 227 1198 372
rect 1209 227 1225 372
rect 1236 227 1252 372
rect 1263 227 1279 372
rect 1290 227 1306 372
rect 1344 227 1360 285
rect 1371 227 1387 285
rect 1399 227 1415 384
rect 1426 227 1442 384
rect 1454 227 1470 368
rect 1481 227 1497 368
rect 1508 227 1524 368
rect 1535 227 1551 368
rect 1563 227 1579 372
rect 1590 227 1606 372
rect 1617 227 1633 372
rect 1644 227 1660 372
rect 1671 227 1687 372
rect 1698 227 1714 372
rect 1725 227 1741 372
rect 1752 227 1768 372
rect 1779 227 1795 372
rect 1846 227 1862 275
rect 1873 227 1889 275
<< metal1 >>
rect 236 454 1831 464
rect 1875 454 1929 464
rect 236 430 1929 440
rect 185 394 1929 419
rect 360 285 376 394
rect 415 384 431 394
rect 470 368 486 394
rect 524 368 540 394
rect 579 372 595 394
rect 633 372 649 394
rect 687 372 703 394
rect 741 372 757 394
rect 795 372 811 394
rect 855 285 871 394
rect 910 384 926 394
rect 965 368 981 394
rect 1019 368 1035 394
rect 1074 372 1090 394
rect 1128 372 1144 394
rect 1182 372 1198 394
rect 1236 372 1252 394
rect 1290 372 1306 394
rect 1344 285 1360 394
rect 1399 384 1415 394
rect 1454 368 1470 394
rect 1508 368 1524 394
rect 1563 372 1579 394
rect 1617 372 1633 394
rect 1671 372 1687 394
rect 1725 372 1741 394
rect 1779 372 1795 394
rect 1855 364 1869 370
rect 1879 275 1889 394
rect 308 198 367 208
rect 393 210 403 227
rect 393 200 422 210
rect 393 187 403 200
rect 448 210 458 227
rect 448 200 477 210
rect 448 187 458 200
rect 503 210 513 227
rect 557 210 567 227
rect 503 200 586 210
rect 503 187 513 200
rect 612 210 622 227
rect 666 210 676 227
rect 720 210 730 227
rect 774 210 784 227
rect 612 200 794 210
rect 612 187 622 200
rect 666 187 676 200
rect 720 187 730 200
rect 774 187 784 200
rect 843 201 862 211
rect 888 210 898 227
rect 888 200 917 210
rect 888 187 898 200
rect 943 210 953 227
rect 943 200 972 210
rect 943 187 953 200
rect 998 210 1008 227
rect 1052 210 1062 227
rect 998 200 1081 210
rect 998 187 1008 200
rect 1107 210 1117 227
rect 1161 210 1171 227
rect 1215 210 1225 227
rect 1269 210 1279 227
rect 1107 200 1295 210
rect 1107 187 1117 200
rect 1161 187 1171 200
rect 1215 187 1225 200
rect 1269 187 1279 200
rect 1336 199 1351 209
rect 1377 210 1387 227
rect 1377 200 1406 210
rect 1377 187 1387 200
rect 1432 210 1442 227
rect 1432 200 1461 210
rect 1432 187 1442 200
rect 1487 210 1497 227
rect 1541 210 1551 227
rect 1487 200 1570 210
rect 1487 187 1497 200
rect 1596 210 1606 227
rect 1650 210 1660 227
rect 1704 210 1714 227
rect 1758 210 1768 227
rect 1596 200 1806 210
rect 1596 187 1606 200
rect 1650 187 1660 200
rect 1704 187 1714 200
rect 1758 187 1768 200
rect 1846 187 1856 227
rect 360 104 376 167
rect 415 104 431 133
rect 470 104 486 114
rect 524 104 540 114
rect 579 104 595 137
rect 633 104 649 137
rect 687 104 703 137
rect 741 104 757 137
rect 795 104 811 137
rect 855 104 871 167
rect 910 104 926 133
rect 965 104 981 114
rect 1019 104 1035 114
rect 1074 104 1090 137
rect 1128 104 1144 137
rect 1182 104 1198 137
rect 1236 104 1252 137
rect 1290 104 1306 137
rect 1344 104 1360 167
rect 1399 104 1415 133
rect 1454 104 1470 114
rect 1508 104 1524 114
rect 1563 104 1579 137
rect 1617 104 1633 137
rect 1671 104 1687 137
rect 1725 104 1741 137
rect 1779 104 1795 137
rect 1873 104 1883 157
rect 360 79 1929 104
rect 808 59 1929 69
rect 284 35 828 45
rect 1309 37 1929 47
rect 260 12 1322 22
rect 1819 15 1929 25
<< m2contact >>
rect 222 453 236 467
rect 1831 451 1845 465
rect 1861 451 1875 465
rect 222 429 236 443
rect 171 394 185 419
rect 1855 370 1869 384
rect 294 196 308 210
rect 794 197 808 211
rect 829 198 843 212
rect 1295 198 1309 212
rect 1322 198 1336 212
rect 1806 198 1820 212
rect 1832 199 1846 213
rect 794 55 808 69
rect 270 33 284 47
rect 828 35 842 49
rect 1295 35 1309 49
rect 246 10 260 24
rect 1322 9 1336 23
rect 1805 13 1819 27
<< metal2 >>
rect 0 419 200 503
rect 223 467 235 503
rect 0 394 171 419
rect 185 394 200 419
rect 0 0 200 394
rect 223 0 235 429
rect 247 24 259 503
rect 271 47 283 503
rect 295 210 307 503
rect 1833 213 1845 451
rect 1861 384 1873 451
rect 1869 370 1873 384
rect 247 0 259 10
rect 271 0 283 33
rect 295 0 307 196
rect 795 69 807 197
rect 830 49 842 198
rect 1296 49 1308 198
rect 1323 23 1335 198
rect 1806 27 1818 198
<< labels >>
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 247 0 259 0 1 Test
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 295 503 307 503 5 nReset
rlabel metal2 271 503 283 503 5 Clock
rlabel metal2 247 503 259 503 5 Test
rlabel metal2 223 503 235 503 5 SDO
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 0 503 200 503 5 Vdd!
rlabel metal2 295 0 307 0 1 nReset
rlabel metal1 1929 430 1929 440 7 SDI
rlabel metal1 1929 454 1929 464 7 nSDO
rlabel metal1 1929 394 1929 419 7 Vdd!
rlabel metal1 1929 79 1929 104 7 GND!
rlabel metal1 1929 15 1929 25 7 TestOut
rlabel metal1 1929 37 1929 47 7 ClockOut
rlabel metal1 1929 59 1929 69 7 nResetOut
<< end >>
