magic
tech c035u
timestamp 1386006598
<< nwell >>
rect 0 402 768 746
<< polysilicon >>
rect 264 681 269 697
rect 399 691 406 719
rect 429 691 436 719
rect 480 704 547 711
rect 76 671 83 679
rect 106 671 113 679
rect 136 671 143 679
rect 180 671 187 679
rect 210 671 217 679
rect 237 671 244 679
rect 264 671 271 681
rect 76 375 83 623
rect 106 553 113 623
rect 136 539 143 623
rect 180 553 187 623
rect 136 523 141 539
rect 106 381 113 505
rect 76 235 83 359
rect 106 335 113 365
rect 136 335 143 523
rect 180 381 187 505
rect 210 381 217 623
rect 237 501 244 623
rect 180 335 187 365
rect 136 319 141 335
rect 106 235 113 305
rect 136 235 143 319
rect 180 235 187 305
rect 210 235 217 365
rect 237 355 244 485
rect 237 235 244 339
rect 264 235 271 623
rect 366 610 373 621
rect 294 583 299 599
rect 294 553 301 583
rect 294 358 301 505
rect 366 388 373 562
rect 399 486 406 643
rect 429 612 436 643
rect 482 612 489 623
rect 523 612 530 645
rect 540 624 547 704
rect 585 691 592 719
rect 643 691 650 719
rect 585 624 592 643
rect 540 617 592 624
rect 585 612 592 617
rect 429 486 436 564
rect 482 486 489 564
rect 523 486 530 564
rect 585 486 592 564
rect 643 532 650 643
rect 711 612 718 675
rect 294 275 301 328
rect 299 259 301 275
rect 366 220 373 372
rect 399 331 406 438
rect 429 402 436 438
rect 482 428 489 438
rect 498 412 510 419
rect 429 395 470 402
rect 463 366 470 395
rect 503 366 510 412
rect 523 410 530 438
rect 585 428 592 438
rect 523 403 551 410
rect 544 366 551 403
rect 585 366 592 412
rect 399 288 406 315
rect 463 288 470 328
rect 76 197 83 205
rect 106 197 113 205
rect 136 197 143 205
rect 180 197 187 205
rect 210 197 217 205
rect 237 197 244 205
rect 264 197 271 205
rect 366 182 373 190
rect 399 161 406 258
rect 463 220 470 258
rect 503 220 510 328
rect 544 220 551 328
rect 585 255 592 328
rect 585 248 599 255
rect 585 225 599 232
rect 585 220 592 225
rect 643 220 650 516
rect 675 486 682 539
rect 675 366 682 438
rect 675 288 682 328
rect 399 110 406 131
rect 463 127 470 190
rect 503 128 510 190
rect 544 161 551 190
rect 585 161 592 190
rect 643 180 650 190
rect 643 142 650 150
rect 675 142 682 258
rect 711 227 718 564
rect 701 220 718 227
rect 708 190 715 195
rect 701 188 715 190
rect 708 180 715 188
rect 708 142 715 150
rect 544 120 551 131
rect 585 120 592 131
<< ndiffusion >>
rect 104 305 106 335
rect 113 305 115 335
rect 178 305 180 335
rect 187 305 189 335
rect 292 328 294 358
rect 301 328 303 358
rect 74 205 76 235
rect 83 205 106 235
rect 113 205 115 235
rect 131 205 136 235
rect 143 205 162 235
rect 178 205 180 235
rect 187 205 210 235
rect 217 205 219 235
rect 235 205 237 235
rect 244 205 264 235
rect 271 205 273 235
rect 458 328 463 366
rect 470 328 503 366
rect 510 328 517 366
rect 533 328 544 366
rect 551 328 585 366
rect 592 328 597 366
rect 394 258 399 288
rect 406 258 463 288
rect 470 258 481 288
rect 364 190 366 220
rect 373 190 378 220
rect 673 258 675 288
rect 682 258 688 288
rect 461 190 463 220
rect 470 190 503 220
rect 510 190 513 220
rect 577 190 585 220
rect 592 190 643 220
rect 650 190 654 220
rect 394 131 399 161
rect 406 131 411 161
rect 542 131 544 161
rect 551 131 585 161
rect 592 131 596 161
rect 705 150 708 180
rect 715 150 718 180
<< pdiffusion >>
rect 74 623 76 671
rect 83 623 88 671
rect 104 623 106 671
rect 113 623 115 671
rect 131 623 136 671
rect 143 623 162 671
rect 178 623 180 671
rect 187 623 189 671
rect 205 623 210 671
rect 217 623 219 671
rect 235 623 237 671
rect 244 623 246 671
rect 262 623 264 671
rect 271 623 273 671
rect 397 643 399 691
rect 406 643 408 691
rect 424 643 429 691
rect 436 643 438 691
rect 104 505 106 553
rect 113 505 115 553
rect 178 505 180 553
rect 187 505 189 553
rect 363 562 366 610
rect 373 562 378 610
rect 292 505 294 553
rect 301 505 303 553
rect 568 643 585 691
rect 592 643 602 691
rect 618 643 643 691
rect 650 643 653 691
rect 427 564 429 612
rect 436 564 464 612
rect 480 564 482 612
rect 489 564 499 612
rect 515 564 523 612
rect 530 564 532 612
rect 548 564 585 612
rect 592 564 594 612
rect 708 564 711 612
rect 718 564 728 612
rect 397 438 399 486
rect 406 438 409 486
rect 425 438 429 486
rect 436 438 438 486
rect 458 438 482 486
rect 489 438 497 486
rect 515 438 523 486
rect 530 438 532 486
rect 548 438 585 486
rect 592 438 595 486
rect 672 438 675 486
rect 682 438 688 486
<< pohmic >>
rect 0 79 54 89
rect 70 79 82 89
rect 98 79 110 89
rect 126 79 138 89
rect 154 79 166 89
rect 182 79 194 89
rect 210 79 222 89
rect 238 79 250 89
rect 266 79 278 89
rect 294 79 306 89
rect 322 79 336 89
rect 0 76 336 79
<< nohmic >>
rect 0 743 336 746
rect 0 736 54 743
rect 70 736 82 743
rect 98 736 110 743
rect 126 736 138 743
rect 154 736 166 743
rect 182 736 194 743
rect 210 736 222 743
rect 238 736 250 743
rect 266 736 278 743
rect 294 736 306 743
rect 322 736 336 743
<< ntransistor >>
rect 106 305 113 335
rect 180 305 187 335
rect 294 328 301 358
rect 76 205 83 235
rect 106 205 113 235
rect 136 205 143 235
rect 180 205 187 235
rect 210 205 217 235
rect 237 205 244 235
rect 264 205 271 235
rect 463 328 470 366
rect 503 328 510 366
rect 544 328 551 366
rect 585 328 592 366
rect 399 258 406 288
rect 463 258 470 288
rect 366 190 373 220
rect 675 258 682 288
rect 463 190 470 220
rect 503 190 510 220
rect 585 190 592 220
rect 643 190 650 220
rect 399 131 406 161
rect 544 131 551 161
rect 585 131 592 161
rect 708 150 715 180
<< ptransistor >>
rect 76 623 83 671
rect 106 623 113 671
rect 136 623 143 671
rect 180 623 187 671
rect 210 623 217 671
rect 237 623 244 671
rect 264 623 271 671
rect 399 643 406 691
rect 429 643 436 691
rect 106 505 113 553
rect 180 505 187 553
rect 366 562 373 610
rect 294 505 301 553
rect 585 643 592 691
rect 643 643 650 691
rect 429 564 436 612
rect 482 564 489 612
rect 523 564 530 612
rect 585 564 592 612
rect 711 564 718 612
rect 399 438 406 486
rect 429 438 436 486
rect 482 438 489 486
rect 523 438 530 486
rect 585 438 592 486
rect 675 438 682 486
<< polycontact >>
rect 269 681 285 697
rect 464 695 480 711
rect 514 645 530 661
rect 141 523 157 539
rect 72 359 88 375
rect 102 365 118 381
rect 228 485 244 501
rect 175 365 191 381
rect 206 365 222 381
rect 141 319 157 335
rect 228 339 244 355
rect 299 583 315 599
rect 702 675 718 691
rect 666 539 682 555
rect 638 516 654 532
rect 357 372 373 388
rect 283 259 299 275
rect 482 412 498 428
rect 585 412 601 428
rect 395 315 411 331
rect 587 232 603 248
rect 666 328 682 366
rect 535 190 551 220
rect 643 150 659 180
rect 692 190 708 220
rect 458 111 474 127
rect 499 111 516 128
<< ndiffcontact >>
rect 88 305 104 335
rect 115 305 131 335
rect 162 305 178 335
rect 189 305 205 335
rect 276 328 292 358
rect 303 328 319 358
rect 58 205 74 235
rect 115 205 131 235
rect 162 205 178 235
rect 219 205 235 235
rect 273 205 289 235
rect 442 328 458 366
rect 517 328 533 366
rect 597 328 613 366
rect 378 258 394 288
rect 481 258 497 288
rect 348 190 364 220
rect 378 190 394 220
rect 657 258 673 288
rect 688 258 704 288
rect 445 190 461 220
rect 513 190 529 220
rect 561 190 577 220
rect 654 190 670 220
rect 378 131 394 161
rect 411 131 427 161
rect 526 131 542 161
rect 596 131 612 161
rect 689 150 705 180
rect 718 150 734 180
<< pdiffcontact >>
rect 57 623 74 671
rect 88 623 104 671
rect 115 623 131 671
rect 162 623 178 671
rect 189 623 205 671
rect 219 623 235 671
rect 246 623 262 671
rect 273 623 289 671
rect 381 643 397 691
rect 408 643 424 691
rect 438 643 454 691
rect 88 505 104 553
rect 115 505 131 553
rect 162 505 178 553
rect 189 505 205 553
rect 347 562 363 610
rect 378 562 394 610
rect 276 505 292 553
rect 303 505 319 553
rect 552 643 568 691
rect 602 643 618 691
rect 653 643 669 691
rect 411 564 427 612
rect 464 564 480 612
rect 499 564 515 612
rect 532 564 548 612
rect 594 564 610 612
rect 692 564 708 612
rect 728 564 744 612
rect 381 438 397 486
rect 409 438 425 486
rect 438 438 458 486
rect 497 438 515 486
rect 532 438 548 486
rect 595 438 611 486
rect 656 438 672 486
rect 688 438 705 486
<< psubstratetap >>
rect 54 79 70 95
rect 82 79 98 95
rect 110 79 126 95
rect 138 79 154 95
rect 166 79 182 95
rect 194 79 210 95
rect 222 79 238 95
rect 250 79 266 95
rect 278 79 294 95
rect 306 79 322 95
rect 552 80 569 97
<< nsubstratetap >>
rect 54 727 70 743
rect 82 727 98 743
rect 110 727 126 743
rect 138 727 154 743
rect 166 727 182 743
rect 194 727 210 743
rect 222 727 238 743
rect 250 727 266 743
rect 278 727 294 743
rect 306 727 322 743
rect 562 727 579 744
<< metal1 >>
rect 0 782 768 792
rect 0 759 222 769
rect 300 759 641 769
rect 657 759 768 769
rect 0 744 768 746
rect 0 743 562 744
rect 0 727 54 743
rect 70 727 82 743
rect 98 727 110 743
rect 126 727 138 743
rect 154 727 166 743
rect 182 727 194 743
rect 210 727 222 743
rect 238 727 250 743
rect 266 727 278 743
rect 294 727 306 743
rect 322 727 562 743
rect 579 727 768 744
rect 0 721 768 727
rect 57 671 74 721
rect 115 671 131 721
rect 141 701 259 711
rect 63 573 74 623
rect 91 613 101 623
rect 141 613 151 701
rect 168 681 232 691
rect 168 671 178 681
rect 222 671 232 681
rect 249 671 259 701
rect 347 634 363 721
rect 381 691 397 721
rect 408 701 464 711
rect 408 691 424 701
rect 602 701 702 711
rect 602 691 618 701
rect 702 691 718 695
rect 347 633 364 634
rect 438 633 454 643
rect 91 603 151 613
rect 192 593 202 623
rect 222 613 232 623
rect 276 613 286 623
rect 222 603 286 613
rect 347 621 454 633
rect 464 645 514 655
rect 347 610 363 621
rect 411 612 427 621
rect 192 583 299 593
rect 63 563 286 573
rect 88 553 98 563
rect 193 553 205 563
rect 157 523 162 539
rect 276 553 286 563
rect 121 495 131 505
rect 121 485 228 495
rect 309 385 319 505
rect 347 511 363 562
rect 464 612 480 645
rect 552 633 568 643
rect 653 633 669 643
rect 728 633 744 721
rect 499 623 744 633
rect 499 612 515 623
rect 594 612 610 623
rect 728 612 744 623
rect 378 549 394 562
rect 464 549 480 564
rect 378 539 480 549
rect 532 554 548 564
rect 532 544 666 554
rect 438 516 612 526
rect 628 516 638 526
rect 692 526 708 564
rect 654 516 708 526
rect 347 501 425 511
rect 409 486 425 501
rect 438 486 458 516
rect 728 506 744 564
rect 497 496 611 506
rect 497 486 515 496
rect 595 486 611 496
rect 656 496 744 506
rect 656 486 672 496
rect 611 438 656 486
rect 381 428 397 438
rect 532 428 548 438
rect 688 428 705 438
rect 381 418 482 428
rect 498 418 548 428
rect 601 418 705 428
rect 396 390 533 402
rect 118 367 120 381
rect 168 365 175 379
rect 309 375 357 385
rect 309 358 319 375
rect 121 345 228 355
rect 121 335 131 345
rect 157 319 162 335
rect 94 295 104 305
rect 195 295 205 305
rect 396 353 409 390
rect 517 366 533 390
rect 348 341 409 353
rect 276 295 286 328
rect 94 285 319 295
rect 61 265 283 275
rect 61 235 71 265
rect 118 245 198 255
rect 118 235 128 245
rect 162 101 178 205
rect 188 195 198 245
rect 222 235 232 265
rect 276 195 286 205
rect 188 185 286 195
rect 309 101 319 285
rect 348 288 364 341
rect 395 314 411 315
rect 613 328 666 366
rect 442 318 458 328
rect 442 308 734 318
rect 348 258 378 288
rect 497 278 657 288
rect 348 220 364 258
rect 378 247 394 258
rect 688 248 704 258
rect 378 235 577 247
rect 561 220 577 235
rect 603 232 704 248
rect 394 190 445 220
rect 529 190 535 220
rect 670 190 692 220
rect 348 161 364 190
rect 718 180 734 308
rect 348 131 378 161
rect 427 151 526 161
rect 659 150 689 180
rect 348 101 366 131
rect 457 111 458 127
rect 596 121 612 131
rect 516 111 612 121
rect 0 97 768 101
rect 0 95 552 97
rect 0 79 54 95
rect 70 79 82 95
rect 98 79 110 95
rect 126 79 138 95
rect 154 79 166 95
rect 182 79 194 95
rect 210 79 222 95
rect 238 79 250 95
rect 266 79 278 95
rect 294 79 306 95
rect 322 80 552 95
rect 569 80 768 97
rect 322 79 768 80
rect 0 76 768 79
rect 0 53 395 63
rect 411 53 768 63
rect 0 30 154 40
rect 168 30 768 40
rect 0 7 441 17
rect 457 7 768 17
<< m2contact >>
rect 222 757 236 771
rect 286 758 300 772
rect 641 756 657 772
rect 285 683 299 697
rect 702 695 718 711
rect 612 516 628 532
rect 120 367 135 381
rect 154 365 168 379
rect 222 367 236 381
rect 72 345 86 359
rect 395 298 411 314
rect 441 111 457 127
rect 395 50 411 66
rect 154 28 168 42
rect 441 3 457 19
<< metal2 >>
rect 72 359 84 799
rect 123 381 135 799
rect 223 743 235 757
rect 222 727 235 743
rect 223 381 235 727
rect 287 697 299 758
rect 614 532 626 799
rect 643 772 655 799
rect 643 711 655 756
rect 643 695 702 711
rect 72 0 84 345
rect 123 0 135 367
rect 155 42 167 365
rect 395 66 411 298
rect 441 19 457 111
rect 614 0 626 516
rect 643 0 655 695
<< labels >>
rlabel metal2 72 799 84 799 5 D
rlabel metal2 123 799 135 799 5 Load
rlabel metal2 72 0 84 0 1 D
rlabel metal2 123 0 135 0 1 Load
rlabel metal2 643 0 655 0 1 Q
rlabel metal2 614 0 626 0 1 nQ
rlabel metal2 643 799 655 799 5 Q
rlabel metal2 614 799 626 799 5 nQ
rlabel metal1 768 7 768 17 7 nReset
rlabel metal1 768 30 768 40 7 Test
rlabel metal1 768 53 768 63 7 Clock
rlabel metal1 768 76 768 101 7 GND!
rlabel metal1 768 759 768 769 7 Q
rlabel metal1 768 782 768 792 7 ScanReturn
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 53 0 63 3 Clock
<< end >>
