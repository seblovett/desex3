magic
tech c035u
timestamp 1385034534
<< nwell >>
rect -10 516 110 729
<< polysilicon >>
rect 53 645 60 653
rect 23 576 30 584
rect 23 518 30 528
rect 23 466 30 502
rect 53 492 60 597
rect 23 428 30 436
rect 53 423 60 476
rect 53 384 60 393
<< ndiffusion >>
rect 21 436 23 466
rect 30 436 32 466
rect 51 393 53 423
rect 60 422 86 423
rect 60 393 70 422
<< pdiffusion >>
rect 48 597 53 645
rect 60 597 70 645
rect 21 528 23 576
rect 30 528 32 576
<< ntransistor >>
rect 23 436 30 466
rect 53 393 60 423
<< ptransistor >>
rect 53 597 60 645
rect 23 528 30 576
<< polycontact >>
rect 22 502 38 518
rect 44 476 60 492
<< ndiffcontact >>
rect 5 436 21 466
rect 32 436 48 466
rect 35 393 51 423
rect 70 393 86 422
<< pdiffcontact >>
rect 32 597 48 645
rect 70 597 86 645
rect 5 528 21 576
rect 32 528 48 576
<< metal1 >>
rect -10 765 110 775
rect -10 742 110 752
rect -10 704 110 729
rect 32 645 48 704
rect 5 597 32 645
rect 5 576 21 597
rect 21 502 22 518
rect 48 492 58 576
rect 70 518 86 597
rect 48 436 58 476
rect 5 423 21 436
rect 5 393 35 423
rect 35 94 51 393
rect 70 422 86 502
rect 70 392 86 393
rect -10 69 110 94
rect -10 46 110 56
rect -10 23 110 33
rect -10 0 110 10
<< m2contact >>
rect 5 502 21 518
rect 70 502 86 518
<< metal2 >>
rect 5 518 21 775
rect 5 0 21 502
rect 70 518 86 775
rect 70 0 86 502
<< labels >>
rlabel metal2 5 0 21 0 1 A
rlabel metal2 5 775 21 775 5 A
rlabel metal2 70 775 86 775 5 Y
rlabel metal2 70 0 86 0 1 Y
rlabel metal1 -10 765 -10 775 4 ScanReturn
rlabel metal1 -10 742 -10 752 3 Scan
rlabel metal1 -10 704 -10 729 3 Vdd!
rlabel metal1 -10 69 -10 94 3 GND!
rlabel metal1 -10 46 -10 56 3 Clock
rlabel metal1 -10 23 -10 33 3 Test
rlabel metal1 -10 0 -10 10 2 nReset
rlabel metal1 110 0 110 10 8 nReset
rlabel metal1 110 23 110 33 7 Test
rlabel metal1 110 46 110 56 7 Clock
rlabel metal1 110 69 110 94 7 GND!
rlabel metal1 110 704 110 729 7 Vdd!
rlabel metal1 110 742 110 752 7 Scan
rlabel metal1 110 765 110 775 6 ScanReturn
<< end >>
