magic
tech c035u
timestamp 1385906671
<< nwell >>
rect 0 302 34 646
<< pohmic >>
rect 0 76 34 92
<< nohmic >>
rect 0 630 34 646
<< metal1 >>
rect 0 682 34 692
rect 0 659 34 669
rect 0 621 34 646
rect 0 95 34 101
rect 0 81 10 95
rect 24 81 34 95
rect 0 76 34 81
rect 0 53 34 63
rect 0 30 34 40
rect 0 7 34 17
<< m2contact >>
rect 10 81 24 95
<< metal2 >>
rect 11 95 23 699
rect 11 0 23 81
<< labels >>
rlabel metal1 34 76 34 101 7 GND!
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 34 53 34 63 7 Clock
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 34 30 34 40 7 Test
rlabel metal1 0 30 0 40 3 Test
rlabel metal2 11 0 23 0 1 GND!
rlabel metal1 0 7 0 17 3 nReset
rlabel metal1 34 7 34 17 7 nReset
rlabel metal1 34 621 34 646 7 Vdd!
rlabel metal1 0 621 0 646 3 Vdd!
rlabel metal1 34 659 34 669 7 Scan
rlabel metal1 0 659 0 669 3 Scan
rlabel metal2 11 699 23 699 5 GND!
rlabel metal1 0 682 0 692 3 ScanReturn
rlabel metal1 34 682 34 692 7 ScanReturn
<< end >>
