magic
tech c035u
timestamp 1385927307
<< nwell >>
rect -7 402 41 746
<< pohmic >>
rect -7 76 41 86
<< nohmic >>
rect -7 736 41 746
<< metal1 >>
rect -7 782 41 792
rect -7 759 41 769
rect -7 740 41 746
rect -7 726 16 740
rect 30 726 41 740
rect -7 721 41 726
rect -7 76 41 101
rect -7 53 41 63
rect -7 30 41 40
rect -7 7 41 17
<< m2contact >>
rect 16 726 30 740
<< metal2 >>
rect 17 740 29 799
rect 17 0 29 726
<< labels >>
rlabel metal1 -7 76 -7 101 3 GND!
rlabel metal1 -7 53 -7 63 3 Clock
rlabel metal1 -7 30 -7 40 3 Test
rlabel metal1 -7 7 -7 17 3 nReset
rlabel metal1 -7 721 -7 746 3 Vdd!
rlabel metal1 -7 759 -7 769 3 Scan
rlabel metal1 -7 782 -7 792 3 ScanReturn
rlabel metal1 41 76 41 101 7 GND!
rlabel metal1 41 53 41 63 7 Clock
rlabel metal1 41 30 41 40 7 Test
rlabel metal1 41 7 41 17 7 nReset
rlabel metal1 41 721 41 746 7 Vdd!
rlabel metal1 41 759 41 769 7 Scan
rlabel metal1 41 782 41 792 7 ScanReturn
rlabel metal2 17 799 29 799 5 Vdd!
rlabel metal2 17 0 29 0 1 Vdd!
<< end >>
