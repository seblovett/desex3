magic
tech c035u
timestamp 1385124685
<< nwell >>
rect 0 521 120 733
<< polysilicon >>
rect 55 569 62 577
rect 55 510 62 521
rect 60 494 62 510
rect 55 481 62 494
rect 55 443 62 451
<< ndiffusion >>
rect 53 451 55 481
rect 62 451 64 481
<< pdiffusion >>
rect 53 521 55 569
rect 62 521 64 569
<< pohmic >>
rect 0 73 6 83
rect 22 73 34 83
rect 50 73 62 83
rect 78 73 90 83
rect 106 73 120 83
<< nohmic >>
rect 0 723 6 733
rect 22 723 34 733
rect 50 723 62 733
rect 78 723 90 733
rect 106 723 120 733
<< ntransistor >>
rect 55 451 62 481
<< ptransistor >>
rect 55 521 62 569
<< polycontact >>
rect 44 494 60 510
<< ndiffcontact >>
rect 37 451 53 481
rect 64 451 80 481
<< pdiffcontact >>
rect 37 521 53 569
rect 64 521 80 569
<< psubstratetap >>
rect 6 73 22 89
rect 34 73 50 89
rect 62 73 78 89
rect 90 73 106 89
<< nsubstratetap >>
rect 6 717 22 733
rect 34 717 50 733
rect 62 717 78 733
rect 90 717 106 733
<< metal1 >>
rect 0 769 120 779
rect 0 746 120 756
rect 0 717 6 733
rect 22 717 34 733
rect 50 717 62 733
rect 78 717 90 733
rect 106 717 120 733
rect 0 708 120 717
rect 37 569 53 708
rect 34 497 44 507
rect 70 508 80 521
rect 70 481 80 494
rect 36 98 52 451
rect 0 89 120 98
rect 0 73 6 89
rect 22 73 34 89
rect 50 73 62 89
rect 78 73 90 89
rect 106 73 120 89
rect 0 50 120 60
rect 0 27 120 37
rect 0 4 120 14
<< m2contact >>
rect 20 495 34 509
rect 70 494 84 508
<< metal2 >>
rect 24 509 36 783
rect 34 495 36 509
rect 72 508 84 783
rect 24 0 36 495
rect 72 0 84 494
<< labels >>
rlabel metal1 0 73 0 98 7 GND!
rlabel metal1 0 50 0 60 7 Clock
rlabel metal1 0 27 0 37 7 Test
rlabel metal1 0 4 0 14 8 nReset
rlabel metal1 0 708 0 733 7 Vdd!
rlabel metal1 0 746 0 756 7 Scan
rlabel metal1 0 769 0 779 6 ScanReturn
rlabel metal2 24 0 36 0 1 A
rlabel metal2 72 0 84 0 1 Y
rlabel metal2 24 783 36 783 5 A
rlabel metal2 72 783 84 783 5 Y
rlabel metal1 120 4 120 14 8 nReset
rlabel metal1 120 27 120 37 7 Test
rlabel metal1 120 50 120 60 7 Clock
rlabel metal1 120 73 120 98 7 GND!
rlabel metal1 120 708 120 733 7 Vdd!
rlabel metal1 120 746 120 756 7 Scan
rlabel metal1 120 769 120 779 6 ScanReturn
<< end >>
