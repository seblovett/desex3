magic
tech c035u
timestamp 1386266982
<< nwell >>
rect 0 401 696 799
<< pwell >>
rect 0 0 696 401
<< polysilicon >>
rect 382 627 389 636
rect 340 558 357 565
rect 307 548 314 556
rect 350 548 357 558
rect 307 490 314 500
rect 55 469 62 477
rect 175 469 182 477
rect 273 469 280 477
rect 350 478 357 500
rect 382 490 389 579
rect 55 391 62 421
rect 175 391 182 421
rect 273 391 280 421
rect 60 375 62 391
rect 180 375 182 391
rect 55 340 62 375
rect 175 340 182 375
rect 273 365 280 375
rect 273 327 280 335
rect 307 330 314 474
rect 55 302 62 310
rect 175 302 182 310
rect 307 304 314 314
rect 350 304 357 328
rect 307 266 314 274
rect 350 264 357 274
rect 382 238 389 474
rect 511 469 518 477
rect 631 469 638 477
rect 511 391 518 421
rect 631 391 638 421
rect 516 375 518 391
rect 636 375 638 391
rect 511 340 518 375
rect 631 340 638 375
rect 511 302 518 310
rect 631 302 638 310
rect 382 200 389 208
<< ndiffusion >>
rect 53 310 55 340
rect 62 310 64 340
rect 173 310 175 340
rect 182 310 184 340
rect 271 335 273 365
rect 280 335 282 365
rect 301 274 307 304
rect 314 274 350 304
rect 357 274 359 304
rect 509 310 511 340
rect 518 310 520 340
rect 629 310 631 340
rect 638 310 640 340
rect 363 208 364 238
rect 380 208 382 238
rect 389 208 391 238
<< pdiffusion >>
rect 380 579 382 627
rect 389 579 391 627
rect 303 500 307 548
rect 314 500 350 548
rect 357 500 359 548
rect 53 421 55 469
rect 62 421 64 469
rect 173 421 175 469
rect 182 421 184 469
rect 271 421 273 469
rect 280 421 282 469
rect 509 421 511 469
rect 518 421 520 469
rect 629 421 631 469
rect 638 421 640 469
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 126 86
rect 142 76 154 86
rect 170 76 182 86
rect 198 76 210 86
rect 226 76 246 86
rect 262 76 274 86
rect 290 76 302 86
rect 318 76 330 86
rect 346 76 358 86
rect 374 76 386 86
rect 402 76 414 86
rect 430 76 462 86
rect 478 76 490 86
rect 506 76 518 86
rect 534 76 546 86
rect 562 76 582 86
rect 598 76 610 86
rect 626 76 638 86
rect 654 76 666 86
rect 682 76 696 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
rect 50 736 62 746
rect 78 736 90 746
rect 106 736 126 746
rect 142 736 154 746
rect 170 736 182 746
rect 198 736 210 746
rect 226 736 246 746
rect 262 736 274 746
rect 290 736 302 746
rect 318 736 330 746
rect 346 736 358 746
rect 374 736 386 746
rect 402 736 414 746
rect 430 736 462 746
rect 478 736 490 746
rect 506 736 518 746
rect 534 736 546 746
rect 562 736 582 746
rect 598 736 610 746
rect 626 736 638 746
rect 654 736 666 746
rect 682 736 696 746
<< ntransistor >>
rect 55 310 62 340
rect 175 310 182 340
rect 273 335 280 365
rect 307 274 314 304
rect 350 274 357 304
rect 511 310 518 340
rect 631 310 638 340
rect 382 208 389 238
<< ptransistor >>
rect 382 579 389 627
rect 307 500 314 548
rect 350 500 357 548
rect 55 421 62 469
rect 175 421 182 469
rect 273 421 280 469
rect 511 421 518 469
rect 631 421 638 469
<< polycontact >>
rect 324 558 340 574
rect 297 474 314 490
rect 44 375 60 391
rect 164 375 180 391
rect 272 375 288 391
rect 298 314 314 330
rect 382 474 398 490
rect 350 248 366 264
rect 500 375 516 391
rect 620 375 636 391
<< ndiffcontact >>
rect 37 310 53 340
rect 64 310 80 340
rect 157 310 173 340
rect 184 310 200 340
rect 255 335 271 365
rect 282 335 298 365
rect 285 274 301 304
rect 359 274 375 304
rect 493 310 509 340
rect 520 310 536 340
rect 613 310 629 340
rect 640 310 656 340
rect 364 208 380 238
rect 391 208 407 238
<< pdiffcontact >>
rect 363 579 380 627
rect 391 579 408 627
rect 285 500 303 548
rect 359 500 375 548
rect 37 421 53 469
rect 64 421 80 469
rect 157 421 173 469
rect 184 421 200 469
rect 255 421 271 469
rect 282 421 298 469
rect 493 421 509 469
rect 520 421 536 469
rect 613 421 629 469
rect 640 421 656 469
<< psubstratetap >>
rect 255 300 271 316
rect 37 281 53 297
rect 157 281 173 297
rect 255 272 271 288
rect 255 244 271 260
rect 493 281 509 297
rect 613 281 629 297
rect 255 216 271 232
rect 255 188 271 204
rect 255 160 271 176
rect 255 132 271 148
rect 255 104 271 120
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 126 76 142 92
rect 154 76 170 92
rect 182 76 198 92
rect 210 76 226 92
rect 246 76 262 92
rect 274 76 290 92
rect 302 76 318 92
rect 330 76 346 92
rect 358 76 374 92
rect 386 76 402 92
rect 414 76 430 92
rect 462 76 478 92
rect 490 76 506 92
rect 518 76 534 92
rect 546 76 562 92
rect 582 76 598 92
rect 610 76 626 92
rect 638 76 654 92
rect 666 76 682 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
rect 62 730 78 746
rect 90 730 106 746
rect 126 730 142 746
rect 154 730 170 746
rect 182 730 198 746
rect 210 730 226 746
rect 246 730 262 746
rect 274 730 290 746
rect 302 730 318 746
rect 330 730 346 746
rect 358 730 374 746
rect 386 730 402 746
rect 414 730 430 746
rect 462 730 478 746
rect 490 730 506 746
rect 518 730 534 746
rect 546 730 562 746
rect 582 730 598 746
rect 610 730 626 746
rect 638 730 654 746
rect 666 730 682 746
<< metal1 >>
rect 85 841 335 851
rect 205 819 263 829
rect 421 818 478 828
rect 494 818 599 828
rect 0 782 696 792
rect 0 759 696 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 62 746
rect 78 730 90 746
rect 106 730 126 746
rect 142 730 154 746
rect 170 730 182 746
rect 198 730 210 746
rect 226 730 246 746
rect 262 730 274 746
rect 290 730 302 746
rect 318 730 330 746
rect 346 730 358 746
rect 374 730 386 746
rect 402 730 414 746
rect 430 730 462 746
rect 478 730 490 746
rect 506 730 518 746
rect 534 730 546 746
rect 562 730 582 746
rect 598 730 610 746
rect 626 730 638 746
rect 654 730 666 746
rect 682 730 696 746
rect 0 721 696 730
rect 37 469 53 721
rect 157 469 173 721
rect 255 469 271 721
rect 285 720 328 721
rect 285 548 303 720
rect 391 627 408 721
rect 350 626 363 627
rect 324 579 363 626
rect 324 574 340 579
rect 282 474 297 490
rect 282 469 298 474
rect 70 389 80 421
rect 190 389 200 421
rect 70 340 80 375
rect 190 340 200 375
rect 255 316 271 335
rect 37 297 53 310
rect 37 101 53 281
rect 157 297 173 310
rect 157 101 173 281
rect 282 314 298 335
rect 255 288 271 300
rect 255 260 271 272
rect 255 232 271 244
rect 255 204 271 216
rect 255 176 271 188
rect 255 148 271 160
rect 255 120 271 132
rect 255 101 271 104
rect 285 101 301 274
rect 324 238 340 558
rect 359 434 372 500
rect 382 473 398 474
rect 493 469 509 721
rect 613 469 629 721
rect 359 417 408 434
rect 359 304 372 417
rect 526 389 536 421
rect 646 389 656 421
rect 526 340 536 375
rect 646 340 656 375
rect 493 297 509 310
rect 366 248 367 264
rect 324 208 364 238
rect 391 101 407 208
rect 493 101 509 281
rect 613 297 629 310
rect 613 101 629 281
rect 0 92 696 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 126 92
rect 142 76 154 92
rect 170 76 182 92
rect 198 76 210 92
rect 226 76 246 92
rect 262 76 274 92
rect 290 76 302 92
rect 318 76 330 92
rect 346 76 358 92
rect 374 76 386 92
rect 402 76 414 92
rect 430 76 462 92
rect 478 76 490 92
rect 506 76 518 92
rect 534 76 546 92
rect 562 76 582 92
rect 598 76 610 92
rect 626 76 638 92
rect 654 76 666 92
rect 682 76 696 92
rect 0 53 696 63
rect 0 30 696 40
rect 0 7 696 17
<< m2contact >>
rect 71 839 85 853
rect 335 839 349 853
rect 191 817 205 831
rect 263 817 277 831
rect 407 815 421 829
rect 478 816 494 830
rect 599 817 613 831
rect 30 376 44 390
rect 70 375 84 389
rect 150 376 164 390
rect 190 375 204 389
rect 256 375 272 391
rect 382 457 398 473
rect 408 417 422 434
rect 486 376 500 390
rect 526 375 540 389
rect 606 376 620 390
rect 646 375 660 389
rect 367 248 383 264
<< metal2 >>
rect 24 390 36 865
rect 24 376 30 390
rect 72 389 84 839
rect 24 0 36 376
rect 72 0 84 375
rect 144 390 156 865
rect 264 831 276 865
rect 336 853 348 865
rect 144 376 150 390
rect 192 389 204 817
rect 264 391 276 817
rect 144 0 156 376
rect 272 375 276 391
rect 192 0 204 375
rect 264 0 276 375
rect 336 473 348 839
rect 408 829 420 865
rect 336 457 382 473
rect 336 264 348 457
rect 408 434 420 815
rect 336 248 367 264
rect 336 0 348 248
rect 408 0 420 417
rect 480 390 492 816
rect 480 376 486 390
rect 528 389 540 799
rect 480 0 492 376
rect 528 0 540 375
rect 600 390 612 817
rect 600 376 606 390
rect 648 389 660 799
rect 600 0 612 376
rect 648 0 660 375
<< labels >>
rlabel metal1 696 721 696 746 7 Vdd!
rlabel metal1 696 759 696 769 7 Scan
rlabel metal1 696 782 696 792 6 ScanReturn
rlabel metal1 696 7 696 17 8 nReset
rlabel metal1 696 30 696 40 7 Test
rlabel metal1 696 53 696 63 7 Clock
rlabel metal1 696 76 696 101 7 GND!
rlabel metal2 24 865 36 865 5 nEnable
rlabel metal2 144 865 156 865 5 nA
rlabel metal2 408 865 420 865 5 Y
rlabel metal2 264 865 276 865 5 A
rlabel metal2 336 865 348 865 5 Enable
<< end >>
