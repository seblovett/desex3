magic
tech c035u
timestamp 1384774380
<< nwell >>
rect 0 320 304 565
<< polysilicon >>
rect 28 490 35 498
rect 58 490 65 540
rect 88 490 95 498
rect 134 490 141 530
rect 218 503 223 519
rect 164 490 171 498
rect 191 490 198 498
rect 218 490 225 503
rect 28 314 35 442
rect 58 372 65 442
rect 88 358 95 442
rect 134 372 141 442
rect 88 342 93 358
rect 28 125 35 298
rect 58 287 65 324
rect 58 221 65 271
rect 88 216 95 342
rect 134 221 141 324
rect 164 267 171 442
rect 191 320 198 442
rect 88 200 93 216
rect 58 125 65 195
rect 88 125 95 200
rect 134 125 141 195
rect 164 125 171 251
rect 191 241 198 304
rect 191 125 198 225
rect 218 125 225 442
rect 262 418 269 425
rect 267 402 269 418
rect 262 372 269 402
rect 262 221 269 324
rect 262 165 269 195
rect 267 149 269 165
rect 28 91 35 99
rect 58 71 65 99
rect 88 91 95 99
rect 134 34 141 99
rect 164 91 171 99
rect 191 91 198 99
rect 218 91 225 99
rect 262 71 269 149
<< ndiffusion >>
rect 56 195 58 221
rect 65 195 67 221
rect 132 195 134 221
rect 141 195 143 221
rect 260 195 262 221
rect 269 195 271 221
rect 26 99 28 125
rect 35 99 58 125
rect 65 99 67 125
rect 83 99 88 125
rect 95 99 116 125
rect 132 99 134 125
rect 141 99 164 125
rect 171 99 173 125
rect 189 99 191 125
rect 198 99 218 125
rect 225 99 227 125
<< pdiffusion >>
rect 26 442 28 490
rect 35 442 40 490
rect 56 442 58 490
rect 65 442 67 490
rect 83 442 88 490
rect 95 442 116 490
rect 132 442 134 490
rect 141 442 143 490
rect 159 442 164 490
rect 171 442 173 490
rect 189 442 191 490
rect 198 442 200 490
rect 216 442 218 490
rect 225 442 227 490
rect 56 324 58 372
rect 65 324 67 372
rect 132 324 134 372
rect 141 324 143 372
rect 260 324 262 372
rect 269 324 271 372
<< ntransistor >>
rect 58 195 65 221
rect 134 195 141 221
rect 262 195 269 221
rect 28 99 35 125
rect 58 99 65 125
rect 88 99 95 125
rect 134 99 141 125
rect 164 99 171 125
rect 191 99 198 125
rect 218 99 225 125
<< ptransistor >>
rect 28 442 35 490
rect 58 442 65 490
rect 88 442 95 490
rect 134 442 141 490
rect 164 442 171 490
rect 191 442 198 490
rect 218 442 225 490
rect 58 324 65 372
rect 134 324 141 372
rect 262 324 269 372
<< polycontact >>
rect 223 503 239 519
rect 93 342 109 358
rect 24 298 40 314
rect 54 271 70 287
rect 182 304 198 320
rect 160 251 176 267
rect 93 200 109 216
rect 182 225 198 241
rect 251 402 267 418
rect 251 149 267 165
rect 126 18 142 34
<< ndiffcontact >>
rect 40 195 56 221
rect 67 195 83 221
rect 116 195 132 221
rect 143 195 159 221
rect 244 195 260 221
rect 271 195 287 221
rect 10 99 26 125
rect 67 99 83 125
rect 116 99 132 125
rect 173 99 189 125
rect 227 99 243 125
<< pdiffcontact >>
rect 9 442 26 490
rect 40 442 56 490
rect 67 442 83 490
rect 116 442 132 490
rect 143 442 159 490
rect 173 442 189 490
rect 200 442 216 490
rect 227 442 243 490
rect 40 324 56 372
rect 67 324 83 372
rect 116 324 132 372
rect 143 324 159 372
rect 244 324 260 372
rect 271 324 287 372
<< psubstratetap >>
rect 7 47 23 63
rect 230 49 246 65
<< nsubstratetap >>
rect 7 543 23 559
rect 230 544 246 560
<< metal1 >>
rect 0 560 304 565
rect 0 559 230 560
rect 0 543 7 559
rect 23 544 230 559
rect 246 544 304 560
rect 23 543 304 544
rect 0 540 304 543
rect 9 490 26 540
rect 67 490 83 540
rect 96 520 213 530
rect 15 392 26 442
rect 43 432 53 442
rect 96 432 106 520
rect 119 500 186 510
rect 119 490 129 500
rect 176 490 186 500
rect 203 490 213 520
rect 239 505 304 515
rect 43 422 106 432
rect 146 412 156 442
rect 176 432 186 442
rect 230 432 240 442
rect 176 422 240 432
rect 146 402 251 412
rect 15 382 254 392
rect 40 372 50 382
rect 147 372 159 382
rect 109 342 116 358
rect 244 372 254 382
rect 73 314 83 324
rect 73 304 182 314
rect 25 288 35 298
rect 70 271 72 285
rect 277 276 287 324
rect 0 251 160 261
rect 277 266 304 276
rect 73 231 182 241
rect 73 221 83 231
rect 277 221 287 266
rect 109 200 116 216
rect 46 185 56 195
rect 149 185 159 195
rect 244 185 254 195
rect 46 175 287 185
rect 13 155 251 165
rect 13 125 23 155
rect 70 135 155 145
rect 70 125 80 135
rect 116 69 132 99
rect 145 89 155 135
rect 176 125 186 155
rect 230 89 240 99
rect 145 79 240 89
rect 277 69 287 175
rect 0 65 304 69
rect 0 63 230 65
rect 0 47 7 63
rect 23 49 230 63
rect 246 49 304 65
rect 23 47 304 49
rect 0 44 304 47
rect 0 24 126 34
<< m2contact >>
rect 23 274 37 288
rect 72 271 87 285
<< metal2 >>
rect 24 288 36 569
rect 75 285 87 569
rect 24 18 36 274
rect 75 18 87 271
<< labels >>
rlabel metal1 304 266 304 276 7 M
rlabel metal1 0 251 0 261 3 SDI
rlabel metal1 0 44 0 69 3 GND!
rlabel metal1 304 44 304 69 7 GND!
rlabel metal2 75 18 87 18 1 Load
rlabel metal2 24 18 36 18 1 D
rlabel metal1 0 24 0 34 3 Test
rlabel metal1 304 540 304 565 1 Vdd!
rlabel metal2 24 569 36 569 5 D
rlabel metal2 75 569 87 569 5 Load
rlabel metal1 304 505 304 515 7 Q
rlabel metal1 0 540 0 565 3 Vdd!
<< end >>
