magic
tech c035u
timestamp 1384961734
<< error_p >>
rect 1919 767 1929 768
rect 1809 25 1819 26
<< nwell >>
rect 1929 743 2073 745
rect 324 533 2073 743
rect 324 505 1820 533
<< polysilicon >>
rect 433 682 440 716
rect 928 682 935 716
rect 1417 682 1424 716
rect 378 583 385 591
rect 488 666 495 674
rect 515 666 522 674
rect 542 666 549 674
rect 597 670 604 678
rect 624 670 631 678
rect 651 670 658 678
rect 678 670 685 678
rect 705 670 712 678
rect 732 670 739 678
rect 759 670 766 678
rect 786 670 793 678
rect 873 583 880 591
rect 983 666 990 674
rect 1010 666 1017 674
rect 1037 666 1044 674
rect 1092 670 1099 678
rect 1119 670 1126 678
rect 1146 670 1153 678
rect 1173 670 1180 678
rect 1200 670 1207 678
rect 1227 670 1234 678
rect 1254 670 1261 678
rect 1281 670 1288 678
rect 1362 583 1369 591
rect 1472 666 1479 674
rect 1499 666 1506 674
rect 1526 666 1533 674
rect 1581 670 1588 678
rect 1608 670 1615 678
rect 1635 670 1642 678
rect 1662 670 1669 678
rect 1689 670 1696 678
rect 1716 670 1723 678
rect 1743 670 1750 678
rect 1770 670 1777 678
rect 1869 646 1871 662
rect 1864 601 1871 646
rect 378 511 385 525
rect 433 511 440 525
rect 488 511 495 525
rect 383 495 385 511
rect 438 495 440 511
rect 493 506 495 511
rect 515 506 522 525
rect 542 506 549 525
rect 597 511 604 525
rect 493 499 549 506
rect 493 495 495 499
rect 378 485 385 495
rect 433 485 440 495
rect 488 485 495 495
rect 515 485 522 499
rect 602 506 604 511
rect 624 506 631 525
rect 651 506 658 525
rect 678 506 685 525
rect 705 506 712 525
rect 732 506 739 525
rect 759 506 766 525
rect 786 508 793 525
rect 873 511 880 525
rect 928 511 935 525
rect 983 511 990 525
rect 784 506 793 508
rect 602 499 793 506
rect 602 495 604 499
rect 597 485 604 495
rect 624 485 631 499
rect 651 485 658 499
rect 678 485 685 499
rect 705 485 712 499
rect 732 485 739 499
rect 759 485 766 499
rect 786 485 793 499
rect 878 495 880 511
rect 933 495 935 511
rect 988 506 990 511
rect 1010 506 1017 525
rect 1037 506 1044 525
rect 1092 511 1099 525
rect 988 499 1044 506
rect 988 495 990 499
rect 873 485 880 495
rect 928 485 935 495
rect 983 485 990 495
rect 1010 485 1017 499
rect 1097 506 1099 511
rect 1119 506 1126 525
rect 1146 506 1153 525
rect 1173 506 1180 525
rect 1200 506 1207 525
rect 1227 506 1234 525
rect 1254 506 1261 525
rect 1281 508 1288 525
rect 1362 511 1369 525
rect 1417 511 1424 525
rect 1472 511 1479 525
rect 1279 506 1288 508
rect 1097 499 1288 506
rect 1097 495 1099 499
rect 1092 485 1099 495
rect 1119 485 1126 499
rect 1146 485 1153 499
rect 1173 485 1180 499
rect 1200 485 1207 499
rect 1227 485 1234 499
rect 1254 485 1261 499
rect 1281 485 1288 499
rect 1367 495 1369 511
rect 1422 495 1424 511
rect 1477 506 1479 511
rect 1499 506 1506 525
rect 1526 506 1533 525
rect 1581 511 1588 525
rect 1477 499 1533 506
rect 1477 495 1479 499
rect 1362 485 1369 495
rect 1417 485 1424 495
rect 1472 485 1479 495
rect 1499 485 1506 499
rect 1586 506 1588 511
rect 1608 506 1615 525
rect 1635 506 1642 525
rect 1662 506 1669 525
rect 1689 506 1696 525
rect 1716 506 1723 525
rect 1743 506 1750 525
rect 1770 508 1777 525
rect 1768 506 1777 508
rect 1586 499 1777 506
rect 1864 505 1871 553
rect 1586 495 1588 499
rect 1581 485 1588 495
rect 1608 485 1615 499
rect 1635 485 1642 499
rect 1662 485 1669 499
rect 1689 485 1696 499
rect 1716 485 1723 499
rect 1743 485 1750 499
rect 1770 485 1777 499
rect 378 457 385 465
rect 433 423 440 431
rect 873 457 880 465
rect 597 427 604 435
rect 624 427 631 435
rect 651 427 658 435
rect 678 427 685 435
rect 705 427 712 435
rect 732 427 739 435
rect 759 427 766 435
rect 786 427 793 435
rect 928 423 935 431
rect 1362 457 1369 465
rect 1092 427 1099 435
rect 1119 427 1126 435
rect 1146 427 1153 435
rect 1173 427 1180 435
rect 1200 427 1207 435
rect 1227 427 1234 435
rect 1254 427 1261 435
rect 1281 427 1288 435
rect 1417 423 1424 431
rect 1864 467 1871 475
rect 1581 427 1588 435
rect 1608 427 1615 435
rect 1635 427 1642 435
rect 1662 427 1669 435
rect 1689 427 1696 435
rect 1716 427 1723 435
rect 1743 427 1750 435
rect 1770 427 1777 435
rect 488 404 495 412
rect 515 404 522 412
rect 983 404 990 412
rect 1010 404 1017 412
rect 1472 404 1479 412
rect 1499 404 1506 412
<< ndiffusion >>
rect 376 465 378 485
rect 385 465 387 485
rect 431 431 433 485
rect 440 431 442 485
rect 486 412 488 485
rect 495 412 497 485
rect 513 412 515 485
rect 522 412 524 485
rect 595 435 597 485
rect 604 435 606 485
rect 622 435 624 485
rect 631 435 633 485
rect 649 435 651 485
rect 658 435 660 485
rect 676 435 678 485
rect 685 435 687 485
rect 703 435 705 485
rect 712 435 714 485
rect 730 435 732 485
rect 739 435 741 485
rect 757 435 759 485
rect 766 435 768 485
rect 784 435 786 485
rect 793 435 795 485
rect 871 465 873 485
rect 880 465 882 485
rect 926 431 928 485
rect 935 431 937 485
rect 981 412 983 485
rect 990 412 992 485
rect 1008 412 1010 485
rect 1017 412 1019 485
rect 1090 435 1092 485
rect 1099 435 1101 485
rect 1117 435 1119 485
rect 1126 435 1128 485
rect 1144 435 1146 485
rect 1153 435 1155 485
rect 1171 435 1173 485
rect 1180 435 1182 485
rect 1198 435 1200 485
rect 1207 435 1209 485
rect 1225 435 1227 485
rect 1234 435 1236 485
rect 1252 435 1254 485
rect 1261 435 1263 485
rect 1279 435 1281 485
rect 1288 435 1290 485
rect 1360 465 1362 485
rect 1369 465 1371 485
rect 1415 431 1417 485
rect 1424 431 1426 485
rect 1470 412 1472 485
rect 1479 412 1481 485
rect 1497 412 1499 485
rect 1506 412 1508 485
rect 1579 435 1581 485
rect 1588 435 1590 485
rect 1606 435 1608 485
rect 1615 435 1617 485
rect 1633 435 1635 485
rect 1642 435 1644 485
rect 1660 435 1662 485
rect 1669 435 1671 485
rect 1687 435 1689 485
rect 1696 435 1698 485
rect 1714 435 1716 485
rect 1723 435 1725 485
rect 1741 435 1743 485
rect 1750 435 1752 485
rect 1768 435 1770 485
rect 1777 435 1779 485
rect 1862 475 1864 505
rect 1871 475 1873 505
<< pdiffusion >>
rect 376 525 378 583
rect 385 525 387 583
rect 431 525 433 682
rect 440 525 442 682
rect 486 525 488 666
rect 495 525 497 666
rect 513 525 515 666
rect 522 525 524 666
rect 540 525 542 666
rect 549 525 551 666
rect 595 525 597 670
rect 604 525 606 670
rect 622 525 624 670
rect 631 525 633 670
rect 649 525 651 670
rect 658 525 660 670
rect 676 525 678 670
rect 685 525 687 670
rect 703 525 705 670
rect 712 525 714 670
rect 730 525 732 670
rect 739 525 741 670
rect 757 525 759 670
rect 766 525 768 670
rect 784 525 786 670
rect 793 525 795 670
rect 871 525 873 583
rect 880 525 882 583
rect 926 525 928 682
rect 935 525 937 682
rect 981 525 983 666
rect 990 525 992 666
rect 1008 525 1010 666
rect 1017 525 1019 666
rect 1035 525 1037 666
rect 1044 525 1046 666
rect 1090 525 1092 670
rect 1099 525 1101 670
rect 1117 525 1119 670
rect 1126 525 1128 670
rect 1144 525 1146 670
rect 1153 525 1155 670
rect 1171 525 1173 670
rect 1180 525 1182 670
rect 1198 525 1200 670
rect 1207 525 1209 670
rect 1225 525 1227 670
rect 1234 525 1236 670
rect 1252 525 1254 670
rect 1261 525 1263 670
rect 1279 525 1281 670
rect 1288 525 1290 670
rect 1360 525 1362 583
rect 1369 525 1371 583
rect 1415 525 1417 682
rect 1424 525 1426 682
rect 1470 525 1472 666
rect 1479 525 1481 666
rect 1497 525 1499 666
rect 1506 525 1508 666
rect 1524 525 1526 666
rect 1533 525 1535 666
rect 1579 525 1581 670
rect 1588 525 1590 670
rect 1606 525 1608 670
rect 1615 525 1617 670
rect 1633 525 1635 670
rect 1642 525 1644 670
rect 1660 525 1662 670
rect 1669 525 1671 670
rect 1687 525 1689 670
rect 1696 525 1698 670
rect 1714 525 1716 670
rect 1723 525 1725 670
rect 1741 525 1743 670
rect 1750 525 1752 670
rect 1768 525 1770 670
rect 1777 525 1779 670
rect 1862 553 1864 601
rect 1871 553 1873 601
<< pohmic >>
rect 376 85 388 95
rect 404 85 416 95
rect 432 85 444 95
rect 460 85 472 95
rect 488 85 500 95
rect 516 85 528 95
rect 544 85 556 95
rect 572 85 584 95
rect 600 85 612 95
rect 628 85 640 95
rect 656 85 668 95
rect 684 85 696 95
rect 712 85 724 95
rect 740 85 752 95
rect 768 85 780 95
rect 796 85 808 95
rect 824 85 836 95
rect 852 85 864 95
rect 880 85 892 95
rect 908 85 920 95
rect 936 85 948 95
rect 964 85 976 95
rect 992 85 1004 95
rect 1020 85 1032 95
rect 1048 85 1060 95
rect 1076 85 1088 95
rect 1104 85 1116 95
rect 1132 85 1144 95
rect 1160 85 1172 95
rect 1188 85 1200 95
rect 1216 85 1228 95
rect 1244 85 1256 95
rect 1272 85 1284 95
rect 1300 85 1312 95
rect 1328 85 1340 95
rect 1356 85 1368 95
rect 1384 85 1396 95
rect 1412 85 1424 95
rect 1440 85 1452 95
rect 1468 85 1480 95
rect 1496 85 1508 95
rect 1524 85 1536 95
rect 1552 85 1564 95
rect 1580 85 1592 95
rect 1608 85 1620 95
rect 1636 85 1648 95
rect 1664 85 1676 95
rect 1692 85 1704 95
rect 1720 85 1732 95
rect 1748 85 1760 95
rect 1776 85 1788 95
rect 1804 85 1816 95
rect 1832 85 1844 95
rect 1860 85 1872 95
rect 1888 85 1900 95
rect 1916 85 1929 95
<< nohmic >>
rect 324 733 334 743
rect 350 733 362 743
rect 378 733 390 743
rect 406 733 418 743
rect 434 733 446 743
rect 462 733 474 743
rect 490 733 502 743
rect 518 733 530 743
rect 546 733 558 743
rect 574 733 586 743
rect 602 733 614 743
rect 630 733 642 743
rect 658 733 670 743
rect 686 733 698 743
rect 714 733 726 743
rect 742 733 754 743
rect 770 733 782 743
rect 798 733 810 743
rect 826 733 838 743
rect 854 733 866 743
rect 882 733 894 743
rect 910 733 922 743
rect 938 733 950 743
rect 966 733 978 743
rect 994 733 1006 743
rect 1022 733 1034 743
rect 1050 733 1062 743
rect 1078 733 1090 743
rect 1106 733 1118 743
rect 1134 733 1146 743
rect 1162 733 1174 743
rect 1190 733 1202 743
rect 1218 733 1230 743
rect 1246 733 1258 743
rect 1274 733 1286 743
rect 1302 733 1314 743
rect 1330 733 1342 743
rect 1358 733 1370 743
rect 1386 733 1398 743
rect 1414 733 1426 743
rect 1442 733 1454 743
rect 1470 733 1482 743
rect 1498 733 1510 743
rect 1526 733 1538 743
rect 1554 733 1566 743
rect 1582 733 1594 743
rect 1610 733 1622 743
rect 1638 733 1650 743
rect 1666 733 1678 743
rect 1694 733 1706 743
rect 1722 733 1734 743
rect 1750 733 1762 743
rect 1778 733 1790 743
rect 1806 733 1818 743
rect 1834 733 1846 743
rect 1862 733 1874 743
rect 1890 733 1902 743
rect 1918 733 1929 743
<< ntransistor >>
rect 378 465 385 485
rect 433 431 440 485
rect 488 412 495 485
rect 515 412 522 485
rect 597 435 604 485
rect 624 435 631 485
rect 651 435 658 485
rect 678 435 685 485
rect 705 435 712 485
rect 732 435 739 485
rect 759 435 766 485
rect 786 435 793 485
rect 873 465 880 485
rect 928 431 935 485
rect 983 412 990 485
rect 1010 412 1017 485
rect 1092 435 1099 485
rect 1119 435 1126 485
rect 1146 435 1153 485
rect 1173 435 1180 485
rect 1200 435 1207 485
rect 1227 435 1234 485
rect 1254 435 1261 485
rect 1281 435 1288 485
rect 1362 465 1369 485
rect 1417 431 1424 485
rect 1472 412 1479 485
rect 1499 412 1506 485
rect 1581 435 1588 485
rect 1608 435 1615 485
rect 1635 435 1642 485
rect 1662 435 1669 485
rect 1689 435 1696 485
rect 1716 435 1723 485
rect 1743 435 1750 485
rect 1770 435 1777 485
rect 1864 475 1871 505
<< ptransistor >>
rect 378 525 385 583
rect 433 525 440 682
rect 488 525 495 666
rect 515 525 522 666
rect 542 525 549 666
rect 597 525 604 670
rect 624 525 631 670
rect 651 525 658 670
rect 678 525 685 670
rect 705 525 712 670
rect 732 525 739 670
rect 759 525 766 670
rect 786 525 793 670
rect 873 525 880 583
rect 928 525 935 682
rect 983 525 990 666
rect 1010 525 1017 666
rect 1037 525 1044 666
rect 1092 525 1099 670
rect 1119 525 1126 670
rect 1146 525 1153 670
rect 1173 525 1180 670
rect 1200 525 1207 670
rect 1227 525 1234 670
rect 1254 525 1261 670
rect 1281 525 1288 670
rect 1362 525 1369 583
rect 1417 525 1424 682
rect 1472 525 1479 666
rect 1499 525 1506 666
rect 1526 525 1533 666
rect 1581 525 1588 670
rect 1608 525 1615 670
rect 1635 525 1642 670
rect 1662 525 1669 670
rect 1689 525 1696 670
rect 1716 525 1723 670
rect 1743 525 1750 670
rect 1770 525 1777 670
rect 1864 553 1871 601
<< polycontact >>
rect 1853 646 1869 662
rect 367 495 383 511
rect 422 495 438 511
rect 477 495 493 511
rect 586 495 602 511
rect 862 495 878 511
rect 917 495 933 511
rect 972 495 988 511
rect 1081 495 1097 511
rect 1351 495 1367 511
rect 1406 495 1422 511
rect 1461 495 1477 511
rect 1570 495 1586 511
<< ndiffcontact >>
rect 360 465 376 485
rect 387 465 403 485
rect 415 431 431 485
rect 442 431 458 485
rect 470 412 486 485
rect 497 412 513 485
rect 524 412 540 485
rect 579 435 595 485
rect 606 435 622 485
rect 633 435 649 485
rect 660 435 676 485
rect 687 435 703 485
rect 714 435 730 485
rect 741 435 757 485
rect 768 435 784 485
rect 795 435 811 485
rect 855 465 871 485
rect 882 465 898 485
rect 910 431 926 485
rect 937 431 953 485
rect 965 412 981 485
rect 992 412 1008 485
rect 1019 412 1035 485
rect 1074 435 1090 485
rect 1101 435 1117 485
rect 1128 435 1144 485
rect 1155 435 1171 485
rect 1182 435 1198 485
rect 1209 435 1225 485
rect 1236 435 1252 485
rect 1263 435 1279 485
rect 1290 435 1306 485
rect 1344 465 1360 485
rect 1371 465 1387 485
rect 1399 431 1415 485
rect 1426 431 1442 485
rect 1454 412 1470 485
rect 1481 412 1497 485
rect 1508 412 1524 485
rect 1563 435 1579 485
rect 1590 435 1606 485
rect 1617 435 1633 485
rect 1644 435 1660 485
rect 1671 435 1687 485
rect 1698 435 1714 485
rect 1725 435 1741 485
rect 1752 435 1768 485
rect 1779 435 1795 485
rect 1846 475 1862 505
rect 1873 475 1889 505
<< pdiffcontact >>
rect 360 525 376 583
rect 387 525 403 583
rect 415 525 431 682
rect 442 525 458 682
rect 470 525 486 666
rect 497 525 513 666
rect 524 525 540 666
rect 551 525 567 666
rect 579 525 595 670
rect 606 525 622 670
rect 633 525 649 670
rect 660 525 676 670
rect 687 525 703 670
rect 714 525 730 670
rect 741 525 757 670
rect 768 525 784 670
rect 795 525 811 670
rect 855 525 871 583
rect 882 525 898 583
rect 910 525 926 682
rect 937 525 953 682
rect 965 525 981 666
rect 992 525 1008 666
rect 1019 525 1035 666
rect 1046 525 1062 666
rect 1074 525 1090 670
rect 1101 525 1117 670
rect 1128 525 1144 670
rect 1155 525 1171 670
rect 1182 525 1198 670
rect 1209 525 1225 670
rect 1236 525 1252 670
rect 1263 525 1279 670
rect 1290 525 1306 670
rect 1344 525 1360 583
rect 1371 525 1387 583
rect 1399 525 1415 682
rect 1426 525 1442 682
rect 1454 525 1470 666
rect 1481 525 1497 666
rect 1508 525 1524 666
rect 1535 525 1551 666
rect 1563 525 1579 670
rect 1590 525 1606 670
rect 1617 525 1633 670
rect 1644 525 1660 670
rect 1671 525 1687 670
rect 1698 525 1714 670
rect 1725 525 1741 670
rect 1752 525 1768 670
rect 1779 525 1795 670
rect 1846 553 1862 601
rect 1873 553 1889 601
<< psubstratetap >>
rect 360 85 376 101
rect 388 85 404 101
rect 416 85 432 101
rect 444 85 460 101
rect 472 85 488 101
rect 500 85 516 101
rect 528 85 544 101
rect 556 85 572 101
rect 584 85 600 101
rect 612 85 628 101
rect 640 85 656 101
rect 668 85 684 101
rect 696 85 712 101
rect 724 85 740 101
rect 752 85 768 101
rect 780 85 796 101
rect 808 85 824 101
rect 836 85 852 101
rect 864 85 880 101
rect 892 85 908 101
rect 920 85 936 101
rect 948 85 964 101
rect 976 85 992 101
rect 1004 85 1020 101
rect 1032 85 1048 101
rect 1060 85 1076 101
rect 1088 85 1104 101
rect 1116 85 1132 101
rect 1144 85 1160 101
rect 1172 85 1188 101
rect 1200 85 1216 101
rect 1228 85 1244 101
rect 1256 85 1272 101
rect 1284 85 1300 101
rect 1312 85 1328 101
rect 1340 85 1356 101
rect 1368 85 1384 101
rect 1396 85 1412 101
rect 1424 85 1440 101
rect 1452 85 1468 101
rect 1480 85 1496 101
rect 1508 85 1524 101
rect 1536 85 1552 101
rect 1564 85 1580 101
rect 1592 85 1608 101
rect 1620 85 1636 101
rect 1648 85 1664 101
rect 1676 85 1692 101
rect 1704 85 1720 101
rect 1732 85 1748 101
rect 1760 85 1776 101
rect 1788 85 1804 101
rect 1816 85 1832 101
rect 1844 85 1860 101
rect 1872 85 1888 101
rect 1900 85 1916 101
<< nsubstratetap >>
rect 334 727 350 743
rect 362 727 378 743
rect 390 727 406 743
rect 418 727 434 743
rect 446 727 462 743
rect 474 727 490 743
rect 502 727 518 743
rect 530 727 546 743
rect 558 727 574 743
rect 586 727 602 743
rect 614 727 630 743
rect 642 727 658 743
rect 670 727 686 743
rect 698 727 714 743
rect 726 727 742 743
rect 754 727 770 743
rect 782 727 798 743
rect 810 727 826 743
rect 838 727 854 743
rect 866 727 882 743
rect 894 727 910 743
rect 922 727 938 743
rect 950 727 966 743
rect 978 727 994 743
rect 1006 727 1022 743
rect 1034 727 1050 743
rect 1062 727 1078 743
rect 1090 727 1106 743
rect 1118 727 1134 743
rect 1146 727 1162 743
rect 1174 727 1190 743
rect 1202 727 1218 743
rect 1230 727 1246 743
rect 1258 727 1274 743
rect 1286 727 1302 743
rect 1314 727 1330 743
rect 1342 727 1358 743
rect 1370 727 1386 743
rect 1398 727 1414 743
rect 1426 727 1442 743
rect 1454 727 1470 743
rect 1482 727 1498 743
rect 1510 727 1526 743
rect 1538 727 1554 743
rect 1566 727 1582 743
rect 1594 727 1610 743
rect 1622 727 1638 743
rect 1650 727 1666 743
rect 1678 727 1694 743
rect 1706 727 1722 743
rect 1734 727 1750 743
rect 1762 727 1778 743
rect 1790 727 1806 743
rect 1818 727 1834 743
rect 1846 727 1862 743
rect 1874 727 1890 743
rect 1902 727 1918 743
<< metal1 >>
rect 236 781 1831 791
rect 1875 781 2073 791
rect 1929 767 2073 768
rect 236 758 2073 767
rect 236 757 1929 758
rect 1929 743 2073 745
rect 185 727 334 743
rect 350 727 362 743
rect 378 727 390 743
rect 406 727 418 743
rect 434 727 446 743
rect 462 727 474 743
rect 490 727 502 743
rect 518 727 530 743
rect 546 727 558 743
rect 574 727 586 743
rect 602 727 614 743
rect 630 727 642 743
rect 658 727 670 743
rect 686 727 698 743
rect 714 727 726 743
rect 742 727 754 743
rect 770 727 782 743
rect 798 727 810 743
rect 826 727 838 743
rect 854 727 866 743
rect 882 727 894 743
rect 910 727 922 743
rect 938 727 950 743
rect 966 727 978 743
rect 994 727 1006 743
rect 1022 727 1034 743
rect 1050 727 1062 743
rect 1078 727 1090 743
rect 1106 727 1118 743
rect 1134 727 1146 743
rect 1162 727 1174 743
rect 1190 727 1202 743
rect 1218 727 1230 743
rect 1246 727 1258 743
rect 1274 727 1286 743
rect 1302 727 1314 743
rect 1330 727 1342 743
rect 1358 727 1370 743
rect 1386 727 1398 743
rect 1414 727 1426 743
rect 1442 727 1454 743
rect 1470 727 1482 743
rect 1498 727 1510 743
rect 1526 727 1538 743
rect 1554 727 1566 743
rect 1582 727 1594 743
rect 1610 727 1622 743
rect 1638 727 1650 743
rect 1666 727 1678 743
rect 1694 727 1706 743
rect 1722 727 1734 743
rect 1750 727 1762 743
rect 1778 727 1790 743
rect 1806 727 1818 743
rect 1834 727 1846 743
rect 1862 727 1874 743
rect 1890 727 1902 743
rect 1918 727 2073 743
rect 185 720 2073 727
rect 185 718 1929 720
rect 360 583 376 718
rect 415 682 431 718
rect 470 666 486 718
rect 524 666 540 718
rect 579 670 595 718
rect 633 670 649 718
rect 687 670 703 718
rect 741 670 757 718
rect 795 670 811 718
rect 855 583 871 718
rect 910 682 926 718
rect 965 666 981 718
rect 1019 666 1035 718
rect 1074 670 1090 718
rect 1128 670 1144 718
rect 1182 670 1198 718
rect 1236 670 1252 718
rect 1290 670 1306 718
rect 1344 583 1360 718
rect 1399 682 1415 718
rect 1454 666 1470 718
rect 1508 666 1524 718
rect 1563 670 1579 718
rect 1617 670 1633 718
rect 1671 670 1687 718
rect 1725 670 1741 718
rect 1779 670 1795 718
rect 1855 662 1869 668
rect 1879 601 1889 718
rect 284 496 367 506
rect 393 508 403 525
rect 393 498 422 508
rect 393 485 403 498
rect 448 508 458 525
rect 448 498 477 508
rect 448 485 458 498
rect 503 508 513 525
rect 557 508 567 525
rect 503 498 586 508
rect 503 485 513 498
rect 612 508 622 525
rect 666 508 676 525
rect 720 508 730 525
rect 774 508 784 525
rect 612 498 794 508
rect 612 485 622 498
rect 666 485 676 498
rect 720 485 730 498
rect 774 485 784 498
rect 843 499 862 509
rect 888 508 898 525
rect 888 498 917 508
rect 888 485 898 498
rect 943 508 953 525
rect 943 498 972 508
rect 943 485 953 498
rect 998 508 1008 525
rect 1052 508 1062 525
rect 998 498 1081 508
rect 998 485 1008 498
rect 1107 508 1117 525
rect 1161 508 1171 525
rect 1215 508 1225 525
rect 1269 508 1279 525
rect 1107 498 1295 508
rect 1107 485 1117 498
rect 1161 485 1171 498
rect 1215 485 1225 498
rect 1269 485 1279 498
rect 1336 497 1351 507
rect 1377 508 1387 525
rect 1377 498 1406 508
rect 1377 485 1387 498
rect 1432 508 1442 525
rect 1432 498 1461 508
rect 1432 485 1442 498
rect 1487 508 1497 525
rect 1541 508 1551 525
rect 1487 498 1570 508
rect 1487 485 1497 498
rect 1596 508 1606 525
rect 1650 508 1660 525
rect 1704 508 1714 525
rect 1758 508 1768 525
rect 1596 498 1806 508
rect 1596 485 1606 498
rect 1650 485 1660 498
rect 1704 485 1714 498
rect 1758 485 1768 498
rect 1846 505 1856 553
rect 360 110 376 465
rect 415 110 431 431
rect 470 110 486 412
rect 524 110 540 412
rect 579 110 595 435
rect 633 110 649 435
rect 687 110 703 435
rect 741 110 757 435
rect 795 110 811 435
rect 855 110 871 465
rect 910 110 926 431
rect 965 110 981 412
rect 1019 110 1035 412
rect 1074 110 1090 435
rect 1128 110 1144 435
rect 1182 110 1198 435
rect 1236 110 1252 435
rect 1290 110 1306 435
rect 1344 110 1360 465
rect 1399 110 1415 431
rect 1454 110 1470 412
rect 1508 110 1524 412
rect 1563 110 1579 435
rect 1617 110 1633 435
rect 1671 110 1687 435
rect 1725 110 1741 435
rect 1779 110 1795 435
rect 1873 110 1883 475
rect 360 101 2073 110
rect 376 85 388 101
rect 404 85 416 101
rect 432 85 444 101
rect 460 85 472 101
rect 488 85 500 101
rect 516 85 528 101
rect 544 85 556 101
rect 572 85 584 101
rect 600 85 612 101
rect 628 85 640 101
rect 656 85 668 101
rect 684 85 696 101
rect 712 85 724 101
rect 740 85 752 101
rect 768 85 780 101
rect 796 85 808 101
rect 824 85 836 101
rect 852 85 864 101
rect 880 85 892 101
rect 908 85 920 101
rect 936 85 948 101
rect 964 85 976 101
rect 992 85 1004 101
rect 1020 85 1032 101
rect 1048 85 1060 101
rect 1076 85 1088 101
rect 1104 85 1116 101
rect 1132 85 1144 101
rect 1160 85 1172 101
rect 1188 85 1200 101
rect 1216 85 1228 101
rect 1244 85 1256 101
rect 1272 85 1284 101
rect 1300 85 1312 101
rect 1328 85 1340 101
rect 1356 85 1368 101
rect 1384 85 1396 101
rect 1412 85 1424 101
rect 1440 85 1452 101
rect 1468 85 1480 101
rect 1496 85 1508 101
rect 1524 85 1536 101
rect 1552 85 1564 101
rect 1580 85 1592 101
rect 1608 85 1620 101
rect 1636 85 1648 101
rect 1664 85 1676 101
rect 1692 85 1704 101
rect 1720 85 1732 101
rect 1748 85 1760 101
rect 1776 85 1788 101
rect 1804 85 1816 101
rect 1832 85 1844 101
rect 1860 85 1872 101
rect 1888 85 1900 101
rect 1916 85 2073 101
rect 808 62 2073 72
rect 260 39 828 49
rect 1309 39 2073 49
rect 308 15 1322 25
rect 1819 16 2073 26
<< m2contact >>
rect 222 779 236 793
rect 1831 778 1845 792
rect 1861 778 1875 792
rect 222 755 236 769
rect 171 718 185 743
rect 1855 668 1869 682
rect 270 494 284 508
rect 794 495 808 509
rect 829 496 843 510
rect 1295 496 1309 510
rect 1322 496 1336 510
rect 1806 496 1820 510
rect 794 61 808 75
rect 246 37 260 51
rect 828 37 842 51
rect 1295 35 1309 49
rect 294 13 308 27
rect 1322 12 1336 26
rect 1805 11 1819 25
<< metal2 >>
rect 0 743 200 827
rect 223 793 235 827
rect 0 718 171 743
rect 185 718 200 743
rect 0 0 200 718
rect 223 0 235 755
rect 247 51 259 827
rect 271 508 283 827
rect 247 0 259 37
rect 271 0 283 494
rect 295 27 307 827
rect 1833 539 1845 778
rect 1861 682 1873 778
rect 1869 668 1873 682
rect 795 75 807 495
rect 830 51 842 496
rect 1296 49 1308 496
rect 1323 26 1335 496
rect 1467 83 1479 103
rect 1502 83 1514 103
rect 295 0 307 13
rect 1806 25 1818 496
<< labels >>
rlabel metal1 1929 85 1929 110 7 GND!
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 295 0 307 0 1 nReset
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 247 0 259 0 1 Test
rlabel metal1 1929 16 1929 26 2 nReset
rlabel metal1 2073 16 2073 26 8 nReset
rlabel metal1 1929 39 1929 49 3 Test
rlabel metal1 2073 39 2073 49 7 Test
rlabel metal1 1929 62 1929 72 3 Clock
rlabel metal1 2073 62 2073 72 7 Clock
rlabel metal1 2073 85 2073 110 7 GND!
rlabel metal1 1929 85 1929 110 3 GND!
rlabel metal1 2073 720 2073 745 7 Vdd!
rlabel metal1 1929 720 1929 745 3 Vdd!
rlabel metal1 2073 758 2073 768 7 Scan
rlabel metal1 1929 758 1929 768 3 Scan
rlabel metal1 1929 781 1929 791 4 ScanReturn
rlabel metal1 2073 781 2073 791 6 ScanReturn
rlabel metal1 1929 62 1929 72 7 ClockOut
rlabel metal1 1929 16 1929 26 7 nResetOut
rlabel metal1 1929 39 1929 49 7 TestOut
rlabel metal2 295 827 307 827 5 nReset
rlabel metal2 271 827 283 827 5 Clock
rlabel metal2 247 827 259 827 5 Test
rlabel metal2 223 827 235 827 5 SDO
rlabel metal2 0 827 200 827 5 Vdd!
rlabel metal1 1929 718 1929 743 7 Vdd!
rlabel metal1 1929 757 1929 767 7 SDI
rlabel metal1 1929 781 1929 791 7 nSDO
<< end >>
