magic
tech c035u
timestamp 1385580953
<< nwell >>
rect 0 460 186 659
<< polysilicon >>
rect 29 604 36 612
rect 59 604 66 612
rect 86 604 93 612
rect 113 604 120 612
rect 144 604 151 612
rect 29 525 36 556
rect 59 512 66 556
rect 29 398 36 477
rect 29 270 36 382
rect 59 270 66 496
rect 86 413 93 556
rect 92 397 93 413
rect 86 270 93 397
rect 113 401 120 556
rect 144 546 151 556
rect 147 530 151 546
rect 113 385 116 401
rect 113 270 120 385
rect 144 316 151 530
rect 146 300 151 316
rect 29 209 36 244
rect 59 205 66 244
rect 86 236 93 244
rect 113 236 120 244
rect 144 209 151 300
rect 29 174 36 183
rect 144 175 151 183
<< ndiffusion >>
rect 27 244 29 270
rect 36 244 38 270
rect 54 244 59 270
rect 66 244 86 270
rect 93 244 95 270
rect 111 244 113 270
rect 120 244 122 270
rect 27 183 29 209
rect 36 183 38 209
rect 142 183 144 209
rect 151 183 153 209
<< pdiffusion >>
rect 27 556 29 604
rect 36 556 38 604
rect 54 556 59 604
rect 66 556 68 604
rect 84 556 86 604
rect 93 556 95 604
rect 111 556 113 604
rect 120 556 123 604
rect 139 556 144 604
rect 151 556 154 604
rect 27 477 29 525
rect 36 477 38 525
<< pohmic >>
rect 0 2 6 9
rect 22 2 34 9
rect 50 2 62 9
rect 78 2 90 9
rect 106 2 118 9
rect 134 2 146 9
rect 162 2 186 9
rect 0 -1 186 2
<< nohmic >>
rect 0 656 186 659
rect 0 649 8 656
rect 24 649 36 656
rect 52 649 64 656
rect 80 649 92 656
rect 108 649 121 656
rect 137 649 149 656
rect 165 649 186 656
<< ntransistor >>
rect 29 244 36 270
rect 59 244 66 270
rect 86 244 93 270
rect 113 244 120 270
rect 29 183 36 209
rect 144 183 151 209
<< ptransistor >>
rect 29 556 36 604
rect 59 556 66 604
rect 86 556 93 604
rect 113 556 120 604
rect 144 556 151 604
rect 29 477 36 525
<< polycontact >>
rect 59 496 75 512
rect 25 382 41 398
rect 76 397 92 413
rect 131 530 147 546
rect 116 385 132 401
rect 130 300 146 316
rect 59 189 75 205
<< ndiffcontact >>
rect 11 244 27 270
rect 38 244 54 270
rect 95 244 111 270
rect 122 244 138 270
rect 11 183 27 209
rect 38 183 54 209
rect 126 183 142 209
rect 153 183 169 209
<< pdiffcontact >>
rect 11 556 27 604
rect 38 556 54 604
rect 68 556 84 604
rect 95 556 111 604
rect 123 556 139 604
rect 154 556 170 604
rect 11 477 27 525
rect 38 477 54 525
<< psubstratetap >>
rect 6 2 22 18
rect 34 2 50 18
rect 62 2 78 18
rect 90 2 106 18
rect 118 2 134 18
rect 146 2 162 18
<< nsubstratetap >>
rect 8 640 24 656
rect 36 640 52 656
rect 64 640 80 656
rect 92 640 108 656
rect 121 640 137 656
rect 149 640 165 656
<< metal1 >>
rect 0 695 186 705
rect 0 672 186 682
rect 0 656 186 659
rect 0 640 8 656
rect 24 640 36 656
rect 52 640 64 656
rect 80 640 92 656
rect 108 640 121 656
rect 137 640 149 656
rect 165 640 186 656
rect 0 634 186 640
rect 11 604 27 634
rect 41 614 108 624
rect 41 604 51 614
rect 98 604 108 614
rect 123 604 139 634
rect 11 525 27 556
rect 71 542 81 556
rect 71 532 131 542
rect 54 496 59 512
rect 157 382 167 556
rect 160 368 167 382
rect 41 303 130 313
rect 41 270 51 303
rect 73 280 135 290
rect 14 234 24 244
rect 73 234 83 280
rect 125 270 135 280
rect 14 224 83 234
rect 95 209 111 244
rect 157 209 167 368
rect 54 189 59 205
rect 95 183 126 209
rect 11 24 27 183
rect 95 24 111 183
rect 0 18 186 24
rect 0 2 6 18
rect 22 2 34 18
rect 50 2 62 18
rect 78 2 90 18
rect 106 2 118 18
rect 134 2 146 18
rect 162 2 186 18
rect 0 -1 186 2
rect 0 -24 186 -14
rect 0 -47 186 -37
rect 0 -70 186 -60
<< m2contact >>
rect 118 401 132 415
rect 41 383 55 397
rect 77 383 91 397
rect 146 368 160 382
<< metal2 >>
rect 48 397 60 709
rect 55 383 60 397
rect 48 -74 60 383
rect 72 397 84 709
rect 120 415 132 709
rect 72 383 77 397
rect 72 -74 84 383
rect 120 -74 132 401
rect 144 382 156 709
rect 144 368 146 382
rect 144 -74 156 368
<< labels >>
rlabel metal1 0 -1 0 24 1 GND!
rlabel metal1 0 -70 0 -60 2 nReset
rlabel metal1 0 -47 0 -37 3 Test
rlabel metal1 0 -24 0 -14 3 Clock
rlabel metal1 0 634 0 659 3 Vdd!
rlabel metal1 0 672 0 682 3 Scan
rlabel metal1 0 695 0 705 4 ScanReturn
rlabel metal2 48 709 60 709 5 S
rlabel metal2 48 -74 60 -74 1 S
rlabel metal2 144 709 156 709 5 Y
rlabel metal2 120 709 132 709 5 I1
rlabel metal2 144 -74 156 -74 1 Y
rlabel metal2 120 -74 132 -74 1 I1
rlabel metal1 186 -1 186 24 7 GND!
rlabel metal1 186 -70 186 -60 8 nReset
rlabel metal1 186 -47 186 -37 7 Test
rlabel metal1 186 -24 186 -14 7 Clock
rlabel metal1 186 634 186 659 7 Vdd!
rlabel metal1 186 695 186 705 6 ScanReturn
rlabel metal1 186 672 186 682 7 Scan
rlabel metal2 72 709 84 709 5 I0
rlabel metal2 72 -74 84 -74 1 I0
<< end >>
