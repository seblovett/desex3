magic
tech c035u
timestamp 1385633707
<< nwell >>
rect 0 402 144 746
<< polysilicon >>
rect 32 450 39 458
rect 59 450 66 458
rect 94 450 101 458
rect 32 372 39 402
rect 36 356 39 372
rect 32 332 39 356
rect 59 372 66 402
rect 94 392 101 402
rect 59 356 67 372
rect 59 332 66 356
rect 94 332 101 376
rect 32 294 39 302
rect 59 294 66 302
rect 94 294 101 302
<< ndiffusion >>
rect 30 302 32 332
rect 39 302 41 332
rect 57 302 59 332
rect 66 302 68 332
rect 92 302 94 332
rect 101 302 103 332
<< pdiffusion >>
rect 30 402 32 450
rect 39 402 59 450
rect 66 402 68 450
rect 92 402 94 450
rect 101 402 103 450
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 144 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
rect 50 736 62 746
rect 78 736 90 746
rect 106 736 144 746
<< ntransistor >>
rect 32 302 39 332
rect 59 302 66 332
rect 94 302 101 332
<< ptransistor >>
rect 32 402 39 450
rect 59 402 66 450
rect 94 402 101 450
<< polycontact >>
rect 20 356 36 372
rect 93 376 109 392
rect 67 356 83 372
<< ndiffcontact >>
rect 6 302 30 332
rect 41 302 57 332
rect 68 302 92 332
rect 103 302 119 332
<< pdiffcontact >>
rect 6 402 30 450
rect 68 402 92 450
rect 103 402 119 450
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
rect 62 730 78 746
rect 90 730 106 746
<< metal1 >>
rect 0 782 144 792
rect 0 759 144 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 62 746
rect 78 730 90 746
rect 106 730 144 746
rect 0 721 144 730
rect 68 450 92 721
rect 6 392 16 402
rect 6 382 93 392
rect 46 332 56 382
rect 119 364 129 450
rect 110 350 129 364
rect 119 302 129 350
rect 6 101 30 302
rect 68 101 92 302
rect 0 92 144 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 144 92
rect 0 53 144 63
rect 0 30 144 40
rect 0 7 144 17
<< m2contact >>
rect 21 342 35 356
rect 67 342 81 356
rect 96 350 110 364
<< metal2 >>
rect 24 356 36 799
rect 35 342 36 356
rect 24 0 36 342
rect 48 356 60 799
rect 96 364 108 799
rect 48 342 67 356
rect 48 0 60 342
rect 96 0 108 350
<< labels >>
rlabel metal1 0 7 0 17 3 nReset
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 144 76 144 101 7 GND!
rlabel metal1 144 53 144 63 7 Clock
rlabel metal1 144 30 144 40 7 Test
rlabel metal1 144 7 144 17 7 nReset
rlabel metal2 24 0 36 0 1 A
rlabel metal2 48 0 60 0 1 B
rlabel metal2 96 0 108 0 1 Y
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 144 721 144 746 1 Vdd!
rlabel metal1 144 759 144 769 1 Scan
rlabel metal1 144 782 144 792 1 ScanReturn
rlabel metal2 24 799 36 799 5 A
rlabel metal2 48 799 60 799 5 B
rlabel metal2 96 799 108 799 5 Y
<< end >>
