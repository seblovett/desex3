magic
tech c035u
timestamp 1384889901
<< nwell >>
rect 0 338 144 550
<< metal1 >>
rect 0 586 144 596
rect 0 563 144 573
rect 0 525 144 550
rect 0 69 144 94
rect 0 46 144 56
rect 0 23 144 33
rect 0 0 144 10
<< labels >>
rlabel metal1 0 0 0 10 2 nReset
rlabel metal1 144 0 144 10 8 nReset
rlabel metal1 0 23 0 33 3 Test
rlabel metal1 144 23 144 33 7 Test
rlabel metal1 0 46 0 56 3 Clock
rlabel metal1 144 46 144 56 7 Clock
rlabel metal1 144 69 144 94 7 GND!
rlabel metal1 0 69 0 94 3 GND!
rlabel metal1 144 525 144 550 7 Vdd!
rlabel metal1 0 525 0 550 3 Vdd!
rlabel metal1 144 563 144 573 7 Scan
rlabel metal1 0 563 0 573 3 Scan
rlabel metal1 0 586 0 596 4 ScanReturn
rlabel metal1 144 586 144 596 6 ScanReturn
<< end >>
