magic
tech c035u
timestamp 1385906433
<< nwell >>
rect 0 302 264 646
<< polysilicon >>
rect 51 597 58 611
rect 24 569 31 577
rect 51 569 58 581
rect 147 569 154 577
rect 177 569 184 577
rect 232 569 239 577
rect 24 491 31 521
rect 51 491 58 521
rect 106 491 113 537
rect 24 249 31 443
rect 24 201 31 231
rect 51 201 58 443
rect 106 201 113 443
rect 147 433 154 521
rect 177 491 184 521
rect 232 461 239 521
rect 238 445 239 461
rect 147 227 154 417
rect 177 279 184 443
rect 24 141 31 171
rect 51 141 58 171
rect 106 161 113 171
rect 147 141 154 211
rect 177 201 184 263
rect 232 217 239 445
rect 177 141 184 171
rect 232 141 239 201
rect 24 103 31 111
rect 51 103 58 111
rect 147 103 154 111
rect 177 103 184 111
rect 232 103 239 111
<< ndiffusion >>
rect 22 171 24 201
rect 31 171 51 201
rect 58 171 60 201
rect 104 171 106 201
rect 113 171 115 201
rect 175 171 177 201
rect 184 171 186 201
rect 22 111 24 141
rect 31 111 33 141
rect 49 111 51 141
rect 58 111 60 141
rect 145 111 147 141
rect 154 111 177 141
rect 184 111 186 141
rect 230 111 232 141
rect 239 111 241 141
<< pdiffusion >>
rect 22 521 24 569
rect 31 521 51 569
rect 58 521 60 569
rect 145 521 147 569
rect 154 521 159 569
rect 175 521 177 569
rect 184 521 186 569
rect 202 521 232 569
rect 239 521 241 569
rect 22 443 24 491
rect 31 443 33 491
rect 49 443 51 491
rect 58 443 60 491
rect 76 443 106 491
rect 113 443 115 491
rect 175 443 177 491
rect 184 443 186 491
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 174 86
rect 190 76 202 86
rect 218 76 230 86
rect 246 76 264 86
<< nohmic >>
rect 0 636 6 646
rect 22 636 34 646
rect 50 636 62 646
rect 78 636 90 646
rect 106 636 118 646
rect 134 636 146 646
rect 162 636 174 646
rect 190 636 202 646
rect 218 636 230 646
rect 246 636 264 646
<< ntransistor >>
rect 24 171 31 201
rect 51 171 58 201
rect 106 171 113 201
rect 177 171 184 201
rect 24 111 31 141
rect 51 111 58 141
rect 147 111 154 141
rect 177 111 184 141
rect 232 111 239 141
<< ptransistor >>
rect 24 521 31 569
rect 51 521 58 569
rect 147 521 154 569
rect 177 521 184 569
rect 232 521 239 569
rect 24 443 31 491
rect 51 443 58 491
rect 106 443 113 491
rect 177 443 184 491
<< polycontact >>
rect 47 581 63 597
rect 101 537 117 553
rect 22 231 40 249
rect 222 445 238 461
rect 138 417 154 433
rect 168 263 184 279
rect 138 211 154 227
rect 101 145 117 161
rect 223 201 239 217
<< ndiffcontact >>
rect 6 171 22 201
rect 60 171 76 201
rect 88 171 104 201
rect 115 171 131 201
rect 159 171 175 201
rect 186 171 202 201
rect 6 111 22 141
rect 33 111 49 141
rect 60 111 76 141
rect 129 111 145 141
rect 186 111 202 141
rect 214 111 230 141
rect 241 111 257 141
<< pdiffcontact >>
rect 6 521 22 569
rect 60 521 76 569
rect 129 521 145 569
rect 159 521 175 569
rect 186 521 202 569
rect 241 521 257 569
rect 6 443 22 491
rect 33 443 49 491
rect 60 443 76 491
rect 115 443 131 491
rect 159 443 175 491
rect 186 443 202 491
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
rect 174 76 190 92
rect 202 76 218 92
rect 230 76 246 92
<< nsubstratetap >>
rect 6 630 22 646
rect 34 630 50 646
rect 62 630 78 646
rect 90 630 106 646
rect 118 630 134 646
rect 146 630 162 646
rect 174 630 190 646
rect 202 630 218 646
rect 230 630 246 646
<< metal1 >>
rect 0 682 264 692
rect 0 659 264 669
rect 0 630 6 646
rect 22 630 34 646
rect 50 630 62 646
rect 78 630 90 646
rect 106 630 118 646
rect 134 630 146 646
rect 162 630 174 646
rect 190 630 202 646
rect 218 630 230 646
rect 246 630 264 646
rect 0 621 264 630
rect 9 569 19 621
rect 132 569 142 621
rect 189 569 199 621
rect 76 540 101 550
rect 9 511 19 521
rect 135 511 145 521
rect 162 511 172 521
rect 9 501 73 511
rect 135 501 152 511
rect 162 501 231 511
rect 9 491 19 501
rect 63 491 73 501
rect 142 491 152 501
rect 142 481 159 491
rect 221 461 231 501
rect 243 485 253 521
rect 221 445 222 461
rect 36 276 46 443
rect 118 430 128 443
rect 192 433 202 443
rect 118 419 138 430
rect 36 266 168 276
rect 63 201 73 266
rect 91 217 138 227
rect 91 201 101 217
rect 192 201 202 227
rect 131 181 159 191
rect 9 141 19 171
rect 36 151 101 161
rect 36 141 46 151
rect 131 141 141 181
rect 222 201 223 217
rect 222 161 232 201
rect 189 151 232 161
rect 189 141 199 151
rect 244 141 254 177
rect 9 101 19 111
rect 63 101 73 111
rect 132 101 142 111
rect 217 101 227 111
rect 0 92 264 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 174 92
rect 190 76 202 92
rect 218 76 230 92
rect 246 76 264 92
rect 0 53 264 63
rect 0 30 264 40
rect 0 7 264 17
<< m2contact >>
rect 47 597 61 611
rect 241 471 255 485
rect 191 419 205 433
rect 24 217 38 231
rect 191 227 205 241
rect 242 177 256 191
<< metal2 >>
rect 24 231 36 699
rect 48 611 60 699
rect 24 0 36 217
rect 48 0 60 597
rect 192 433 204 699
rect 240 485 252 699
rect 240 471 241 485
rect 192 241 204 419
rect 192 0 204 227
rect 240 191 252 471
rect 240 177 242 191
rect 240 0 252 177
<< labels >>
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 264 76 264 101 7 GND!
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 264 53 264 63 7 Clock
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 264 30 264 40 7 Test
rlabel metal2 24 0 36 0 1 A
rlabel metal2 48 0 60 0 1 B
rlabel metal2 192 0 204 0 1 C
rlabel metal2 240 0 252 0 1 S
rlabel metal1 0 7 0 17 3 nReset
rlabel metal1 264 7 264 17 7 nReset
rlabel metal1 0 621 0 646 3 Vdd!
rlabel metal1 264 621 264 646 7 Vdd!
rlabel metal1 0 659 0 669 3 Scan
rlabel metal1 264 659 264 669 7 Scan
rlabel metal1 0 682 0 692 3 ScanReturn
rlabel metal1 264 682 264 692 7 ScanReturn
rlabel metal2 240 699 252 699 5 S
rlabel metal2 192 699 204 699 5 C
rlabel metal2 48 699 60 699 5 B
rlabel metal2 24 699 36 699 5 A
<< end >>
