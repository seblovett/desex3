magic
tech c035u
timestamp 1386241447
<< nwell >>
rect 0 401 720 799
<< pwell >>
rect 0 0 720 401
<< polysilicon >>
rect 216 681 221 697
rect 355 691 362 719
rect 385 691 392 719
rect 436 704 503 711
rect 28 671 35 679
rect 58 671 65 679
rect 88 671 95 679
rect 132 671 139 679
rect 162 671 169 679
rect 189 671 196 679
rect 216 671 223 681
rect 28 375 35 623
rect 58 553 65 623
rect 88 539 95 623
rect 132 553 139 623
rect 88 523 93 539
rect 58 381 65 505
rect 28 235 35 359
rect 58 335 65 365
rect 88 335 95 523
rect 132 381 139 505
rect 162 381 169 623
rect 189 501 196 623
rect 132 335 139 365
rect 88 319 93 335
rect 58 235 65 305
rect 88 235 95 319
rect 132 235 139 305
rect 162 235 169 365
rect 189 355 196 485
rect 189 235 196 339
rect 216 235 223 623
rect 322 610 329 621
rect 246 583 251 599
rect 246 553 253 583
rect 246 358 253 505
rect 322 388 329 562
rect 355 486 362 643
rect 385 612 392 643
rect 438 612 445 623
rect 479 612 486 645
rect 496 624 503 704
rect 541 691 548 719
rect 599 691 606 719
rect 541 624 548 643
rect 496 617 548 624
rect 541 612 548 617
rect 385 486 392 564
rect 438 486 445 564
rect 479 486 486 564
rect 541 486 548 564
rect 599 532 606 643
rect 667 612 674 675
rect 246 275 253 328
rect 251 259 253 275
rect 322 225 329 372
rect 355 331 362 438
rect 385 402 392 438
rect 438 428 445 438
rect 454 412 466 419
rect 385 395 426 402
rect 419 358 426 395
rect 459 358 466 412
rect 479 410 486 438
rect 541 428 548 438
rect 479 403 507 410
rect 500 358 507 403
rect 541 358 548 412
rect 355 288 362 315
rect 419 288 426 328
rect 28 197 35 205
rect 58 197 65 205
rect 88 197 95 205
rect 132 197 139 205
rect 162 197 169 205
rect 189 197 196 205
rect 216 197 223 205
rect 322 187 329 195
rect 355 161 362 258
rect 419 225 426 258
rect 459 225 466 328
rect 500 225 507 328
rect 541 255 548 328
rect 541 248 555 255
rect 541 225 555 232
rect 541 220 548 225
rect 599 220 606 516
rect 631 486 638 539
rect 631 358 638 438
rect 631 288 638 328
rect 355 110 362 131
rect 419 127 426 195
rect 459 128 466 195
rect 500 161 507 195
rect 541 161 548 190
rect 599 180 606 190
rect 599 142 606 150
rect 631 142 638 258
rect 667 227 674 564
rect 657 220 674 227
rect 664 190 671 195
rect 657 188 671 190
rect 664 180 671 188
rect 664 142 671 150
rect 500 120 507 131
rect 541 120 548 131
<< ndiffusion >>
rect 56 305 58 335
rect 65 305 67 335
rect 130 305 132 335
rect 139 305 141 335
rect 244 328 246 358
rect 253 328 255 358
rect 26 205 28 235
rect 35 205 58 235
rect 65 205 67 235
rect 83 205 88 235
rect 95 205 114 235
rect 130 205 132 235
rect 139 205 162 235
rect 169 205 171 235
rect 187 205 189 235
rect 196 205 216 235
rect 223 205 225 235
rect 414 328 419 358
rect 426 328 459 358
rect 466 328 473 358
rect 489 328 500 358
rect 507 328 541 358
rect 548 328 553 358
rect 350 258 355 288
rect 362 258 419 288
rect 426 258 437 288
rect 320 195 322 225
rect 329 195 334 225
rect 417 195 419 225
rect 426 195 459 225
rect 466 195 469 225
rect 629 258 631 288
rect 638 258 644 288
rect 350 131 355 161
rect 362 131 367 161
rect 533 190 541 220
rect 548 190 599 220
rect 606 190 610 220
rect 498 131 500 161
rect 507 131 541 161
rect 548 131 552 161
rect 661 150 664 180
rect 671 150 674 180
<< pdiffusion >>
rect 26 623 28 671
rect 35 623 40 671
rect 56 623 58 671
rect 65 623 67 671
rect 83 623 88 671
rect 95 623 114 671
rect 130 623 132 671
rect 139 623 141 671
rect 157 623 162 671
rect 169 623 171 671
rect 187 623 189 671
rect 196 623 198 671
rect 214 623 216 671
rect 223 623 225 671
rect 353 643 355 691
rect 362 643 364 691
rect 380 643 385 691
rect 392 643 394 691
rect 56 505 58 553
rect 65 505 67 553
rect 130 505 132 553
rect 139 505 141 553
rect 319 562 322 610
rect 329 562 334 610
rect 244 505 246 553
rect 253 505 255 553
rect 524 643 541 691
rect 548 643 558 691
rect 574 643 599 691
rect 606 643 609 691
rect 383 564 385 612
rect 392 564 420 612
rect 436 564 438 612
rect 445 564 455 612
rect 471 564 479 612
rect 486 564 488 612
rect 504 564 541 612
rect 548 564 550 612
rect 664 564 667 612
rect 674 564 684 612
rect 353 438 355 486
rect 362 438 365 486
rect 381 438 385 486
rect 392 438 394 486
rect 414 438 438 486
rect 445 438 453 486
rect 471 438 479 486
rect 486 438 488 486
rect 504 438 541 486
rect 548 438 551 486
rect 628 438 631 486
rect 638 438 644 486
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 174 86
rect 190 79 202 86
rect 218 79 230 86
rect 246 79 258 86
rect 274 79 298 86
rect 0 76 298 79
rect 314 76 326 86
rect 342 76 354 86
rect 370 76 382 86
rect 398 76 410 86
rect 426 76 438 86
rect 454 76 466 86
rect 482 76 494 86
rect 510 76 522 86
rect 539 76 551 86
rect 567 76 579 86
rect 595 76 607 86
rect 623 76 635 86
rect 652 76 664 86
rect 681 76 693 86
rect 710 76 720 86
<< nohmic >>
rect 0 743 298 746
rect 0 736 6 743
rect 22 736 34 743
rect 50 736 62 743
rect 78 736 90 743
rect 106 736 118 743
rect 134 736 146 743
rect 162 736 174 743
rect 190 736 202 743
rect 218 736 230 743
rect 246 736 258 743
rect 274 736 298 743
rect 314 736 326 746
rect 342 736 354 746
rect 370 736 382 746
rect 398 736 410 746
rect 426 736 438 746
rect 454 736 466 746
rect 482 736 494 746
rect 510 736 522 746
rect 538 736 550 746
rect 566 736 578 746
rect 594 736 606 746
rect 622 736 634 746
rect 650 736 662 746
rect 678 736 690 746
rect 706 736 720 746
<< ntransistor >>
rect 58 305 65 335
rect 132 305 139 335
rect 246 328 253 358
rect 28 205 35 235
rect 58 205 65 235
rect 88 205 95 235
rect 132 205 139 235
rect 162 205 169 235
rect 189 205 196 235
rect 216 205 223 235
rect 419 328 426 358
rect 459 328 466 358
rect 500 328 507 358
rect 541 328 548 358
rect 355 258 362 288
rect 419 258 426 288
rect 322 195 329 225
rect 419 195 426 225
rect 459 195 466 225
rect 631 258 638 288
rect 355 131 362 161
rect 541 190 548 220
rect 599 190 606 220
rect 500 131 507 161
rect 541 131 548 161
rect 664 150 671 180
<< ptransistor >>
rect 28 623 35 671
rect 58 623 65 671
rect 88 623 95 671
rect 132 623 139 671
rect 162 623 169 671
rect 189 623 196 671
rect 216 623 223 671
rect 355 643 362 691
rect 385 643 392 691
rect 58 505 65 553
rect 132 505 139 553
rect 322 562 329 610
rect 246 505 253 553
rect 541 643 548 691
rect 599 643 606 691
rect 385 564 392 612
rect 438 564 445 612
rect 479 564 486 612
rect 541 564 548 612
rect 667 564 674 612
rect 355 438 362 486
rect 385 438 392 486
rect 438 438 445 486
rect 479 438 486 486
rect 541 438 548 486
rect 631 438 638 486
<< polycontact >>
rect 221 681 237 697
rect 420 695 436 711
rect 470 645 486 661
rect 93 523 109 539
rect 24 359 40 375
rect 54 365 70 381
rect 180 485 196 501
rect 127 365 143 381
rect 158 365 174 381
rect 93 319 109 335
rect 180 339 196 355
rect 251 583 267 599
rect 658 675 674 691
rect 622 539 638 555
rect 594 516 610 532
rect 313 372 329 388
rect 235 259 251 275
rect 438 412 454 428
rect 541 412 557 428
rect 351 315 367 331
rect 543 232 559 248
rect 491 195 507 225
rect 622 328 638 358
rect 599 150 615 180
rect 648 190 664 220
rect 414 111 430 127
rect 455 111 472 128
<< ndiffcontact >>
rect 40 305 56 335
rect 67 305 83 335
rect 114 305 130 335
rect 141 305 157 335
rect 228 328 244 358
rect 255 328 271 358
rect 10 205 26 235
rect 67 205 83 235
rect 114 205 130 235
rect 171 205 187 235
rect 225 205 241 235
rect 398 328 414 358
rect 473 328 489 358
rect 553 328 569 358
rect 334 258 350 288
rect 437 258 453 288
rect 304 195 320 225
rect 334 195 350 225
rect 401 195 417 225
rect 469 195 485 225
rect 613 258 629 288
rect 644 258 660 288
rect 334 131 350 161
rect 367 131 383 161
rect 517 190 533 220
rect 610 190 626 220
rect 482 131 498 161
rect 552 131 568 161
rect 645 150 661 180
rect 674 150 690 180
<< pdiffcontact >>
rect 9 623 26 671
rect 40 623 56 671
rect 67 623 83 671
rect 114 623 130 671
rect 141 623 157 671
rect 171 623 187 671
rect 198 623 214 671
rect 225 623 241 671
rect 337 643 353 691
rect 364 643 380 691
rect 394 643 410 691
rect 40 505 56 553
rect 67 505 83 553
rect 114 505 130 553
rect 141 505 157 553
rect 303 562 319 610
rect 334 562 350 610
rect 228 505 244 553
rect 255 505 271 553
rect 508 643 524 691
rect 558 643 574 691
rect 609 643 625 691
rect 367 564 383 612
rect 420 564 436 612
rect 455 564 471 612
rect 488 564 504 612
rect 550 564 566 612
rect 648 564 664 612
rect 684 564 700 612
rect 337 438 353 486
rect 365 438 381 486
rect 394 438 414 486
rect 453 438 471 486
rect 488 438 504 486
rect 551 438 567 486
rect 612 438 628 486
rect 644 438 661 486
<< psubstratetap >>
rect 301 337 317 353
rect 114 175 130 192
rect 304 166 320 182
rect 6 79 22 96
rect 34 79 50 96
rect 62 79 78 96
rect 90 79 106 96
rect 118 79 134 96
rect 146 79 162 96
rect 174 79 190 96
rect 202 79 218 96
rect 230 79 246 96
rect 258 79 274 96
rect 298 76 314 92
rect 326 76 342 92
rect 354 76 370 92
rect 382 76 398 92
rect 410 76 426 92
rect 438 76 454 92
rect 466 76 482 92
rect 494 76 510 92
rect 522 76 539 92
rect 551 76 567 92
rect 579 76 595 92
rect 607 76 623 92
rect 635 76 652 92
rect 664 76 681 92
rect 693 76 710 92
<< nsubstratetap >>
rect 6 727 22 743
rect 34 727 50 743
rect 62 727 78 743
rect 90 727 106 743
rect 118 727 134 743
rect 146 727 162 743
rect 174 727 190 743
rect 202 727 218 743
rect 230 727 246 743
rect 258 727 274 743
rect 298 730 314 746
rect 326 730 342 746
rect 354 730 370 746
rect 382 730 398 746
rect 410 730 426 746
rect 438 730 454 746
rect 466 730 482 746
rect 494 730 510 746
rect 522 730 538 746
rect 550 730 566 746
rect 578 730 594 746
rect 606 730 622 746
rect 634 730 650 746
rect 662 730 678 746
rect 690 730 706 746
<< metal1 >>
rect 0 782 720 792
rect 0 759 174 769
rect 252 759 598 769
rect 614 759 720 769
rect 0 743 298 746
rect 0 727 6 743
rect 22 727 34 743
rect 50 727 62 743
rect 78 727 90 743
rect 106 727 118 743
rect 134 727 146 743
rect 162 727 174 743
rect 190 727 202 743
rect 218 727 230 743
rect 246 727 258 743
rect 274 730 298 743
rect 314 730 326 746
rect 342 730 354 746
rect 370 730 382 746
rect 398 730 410 746
rect 426 730 438 746
rect 454 730 466 746
rect 482 730 494 746
rect 510 730 522 746
rect 538 730 550 746
rect 566 730 578 746
rect 594 730 606 746
rect 622 730 634 746
rect 650 730 662 746
rect 678 730 690 746
rect 706 730 720 746
rect 274 727 720 730
rect 0 721 720 727
rect 9 671 26 721
rect 67 671 83 721
rect 93 701 211 711
rect 15 573 26 623
rect 43 613 53 623
rect 93 613 103 701
rect 120 681 184 691
rect 120 671 130 681
rect 174 671 184 681
rect 201 671 211 701
rect 303 634 319 721
rect 337 691 353 721
rect 364 701 420 711
rect 364 691 380 701
rect 558 701 658 711
rect 558 691 574 701
rect 658 691 674 695
rect 303 633 320 634
rect 394 633 410 643
rect 43 603 103 613
rect 144 593 154 623
rect 174 613 184 623
rect 228 613 238 623
rect 174 603 238 613
rect 303 621 410 633
rect 420 645 470 655
rect 303 610 319 621
rect 367 612 383 621
rect 144 583 251 593
rect 15 563 238 573
rect 40 553 50 563
rect 145 553 157 563
rect 109 523 114 539
rect 228 553 238 563
rect 73 495 83 505
rect 73 485 180 495
rect 261 385 271 505
rect 303 511 319 562
rect 420 612 436 645
rect 508 633 524 643
rect 609 633 625 643
rect 684 633 700 721
rect 455 623 700 633
rect 455 612 471 623
rect 550 612 566 623
rect 684 612 700 623
rect 334 549 350 562
rect 420 549 436 564
rect 334 539 436 549
rect 488 554 504 564
rect 488 544 622 554
rect 394 516 550 526
rect 566 516 594 526
rect 648 526 664 564
rect 610 516 664 526
rect 303 501 381 511
rect 365 486 381 501
rect 394 486 414 516
rect 684 506 700 564
rect 453 496 567 506
rect 453 486 471 496
rect 551 486 567 496
rect 612 496 700 506
rect 612 486 628 496
rect 567 438 612 486
rect 337 428 353 438
rect 488 428 504 438
rect 644 428 661 438
rect 337 418 438 428
rect 454 418 504 428
rect 557 418 661 428
rect 352 390 489 402
rect 120 365 127 379
rect 261 375 313 385
rect 261 358 271 375
rect 73 345 180 355
rect 73 335 83 345
rect 109 319 114 335
rect 46 295 56 305
rect 147 295 157 305
rect 352 353 365 390
rect 473 358 489 390
rect 317 341 365 353
rect 317 337 320 341
rect 228 295 238 328
rect 46 285 271 295
rect 13 265 235 275
rect 13 235 23 265
rect 70 245 150 255
rect 70 235 80 245
rect 114 192 130 205
rect 140 195 150 245
rect 174 235 184 265
rect 228 195 238 205
rect 140 185 238 195
rect 114 101 130 175
rect 261 101 271 285
rect 304 288 320 337
rect 351 314 367 315
rect 569 328 622 358
rect 398 318 414 328
rect 398 308 690 318
rect 304 258 334 288
rect 453 278 613 288
rect 304 225 320 258
rect 334 247 350 258
rect 644 248 660 258
rect 334 235 533 247
rect 350 195 401 225
rect 485 195 491 225
rect 517 220 533 235
rect 559 232 660 248
rect 304 182 320 195
rect 626 190 648 220
rect 674 180 690 308
rect 304 161 320 166
rect 304 131 334 161
rect 383 151 482 161
rect 615 150 645 180
rect 304 101 322 131
rect 413 111 414 127
rect 552 121 568 131
rect 472 111 568 121
rect 0 96 720 101
rect 0 79 6 96
rect 22 79 34 96
rect 50 79 62 96
rect 78 79 90 96
rect 106 79 118 96
rect 134 79 146 96
rect 162 79 174 96
rect 190 79 202 96
rect 218 79 230 96
rect 246 79 258 96
rect 274 92 720 96
rect 274 79 298 92
rect 0 76 298 79
rect 314 76 326 92
rect 342 76 354 92
rect 370 76 382 92
rect 398 76 410 92
rect 426 76 438 92
rect 454 76 466 92
rect 482 76 494 92
rect 510 76 522 92
rect 539 76 551 92
rect 567 76 579 92
rect 595 76 607 92
rect 623 76 635 92
rect 652 76 664 92
rect 681 76 693 92
rect 710 76 720 92
rect 0 53 351 63
rect 367 53 720 63
rect 0 30 106 40
rect 120 30 720 40
rect 0 7 397 17
rect 413 7 720 17
<< m2contact >>
rect 174 757 188 771
rect 238 758 252 772
rect 598 756 614 772
rect 237 683 251 697
rect 658 695 674 711
rect 550 516 566 532
rect 70 367 85 381
rect 106 365 120 379
rect 174 367 188 381
rect 24 345 38 359
rect 351 298 367 314
rect 397 111 413 127
rect 351 50 367 66
rect 106 28 120 42
rect 397 4 413 20
<< metal2 >>
rect 24 359 36 799
rect 72 381 84 799
rect 175 743 187 757
rect 174 727 187 743
rect 175 381 187 727
rect 239 697 251 758
rect 552 532 564 799
rect 600 772 612 799
rect 600 711 612 756
rect 600 695 658 711
rect 24 0 36 345
rect 72 0 84 367
rect 107 42 119 365
rect 351 66 367 298
rect 397 20 413 111
rect 552 0 564 516
rect 600 0 612 695
<< labels >>
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal2 24 799 36 799 5 D
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 53 0 63 3 Clock
rlabel metal2 24 0 36 0 1 D
rlabel metal2 72 0 84 0 1 Load
rlabel metal2 72 799 84 799 5 Load
rlabel metal1 720 782 720 792 7 ScanReturn
rlabel metal1 720 759 720 769 7 Q
rlabel metal1 720 76 720 101 7 GND!
rlabel metal1 720 53 720 63 7 Clock
rlabel metal1 720 30 720 40 7 Test
rlabel metal1 720 7 720 17 7 nReset
rlabel metal1 720 721 720 746 7 Vdd!
rlabel metal2 552 0 564 0 1 nQ
rlabel metal2 600 0 612 0 1 Q
rlabel metal2 600 799 612 799 5 Q
rlabel metal2 552 799 564 799 5 nQ
<< end >>
