magic
tech c035u
timestamp 1385030757
<< nwell >>
rect 16 657 423 733
rect 16 422 422 657
rect 16 421 58 422
<< polysilicon >>
rect 77 678 84 706
rect 107 678 114 706
rect 158 691 225 698
rect 44 597 51 608
rect 44 388 51 549
rect 77 473 84 630
rect 107 599 114 630
rect 160 599 167 610
rect 201 599 208 632
rect 218 611 225 691
rect 263 678 270 706
rect 321 678 328 706
rect 263 611 270 630
rect 218 604 270 611
rect 263 599 270 604
rect 107 473 114 551
rect 160 473 167 551
rect 201 473 208 551
rect 263 473 270 551
rect 321 519 328 630
rect 389 599 396 662
rect 44 217 51 372
rect 77 328 84 425
rect 107 389 114 425
rect 160 415 167 425
rect 176 399 188 406
rect 107 382 148 389
rect 141 363 148 382
rect 181 363 188 399
rect 201 397 208 425
rect 263 415 270 425
rect 201 390 229 397
rect 222 363 229 390
rect 263 363 270 399
rect 77 285 84 312
rect 141 285 148 325
rect 44 179 51 187
rect 77 158 84 255
rect 141 217 148 255
rect 181 217 188 325
rect 222 217 229 325
rect 263 252 270 325
rect 263 245 277 252
rect 263 222 277 229
rect 263 217 270 222
rect 321 217 328 503
rect 353 473 360 526
rect 353 363 360 425
rect 353 285 360 325
rect 77 107 84 128
rect 141 124 148 187
rect 181 125 188 187
rect 222 158 229 187
rect 263 158 270 187
rect 321 177 328 187
rect 321 139 328 147
rect 353 139 360 255
rect 389 224 396 551
rect 379 217 396 224
rect 386 187 393 192
rect 379 185 393 187
rect 386 177 393 185
rect 386 139 393 147
rect 222 117 229 128
rect 263 117 270 128
<< ndiffusion >>
rect 136 325 141 363
rect 148 325 181 363
rect 188 325 195 363
rect 211 325 222 363
rect 229 325 263 363
rect 270 325 275 363
rect 72 255 77 285
rect 84 255 141 285
rect 148 255 159 285
rect 42 187 44 217
rect 51 187 56 217
rect 351 255 353 285
rect 360 255 366 285
rect 139 187 141 217
rect 148 187 181 217
rect 188 187 191 217
rect 255 187 263 217
rect 270 187 321 217
rect 328 187 332 217
rect 72 128 77 158
rect 84 128 89 158
rect 220 128 222 158
rect 229 128 263 158
rect 270 128 274 158
rect 383 147 386 177
rect 393 147 396 177
<< pdiffusion >>
rect 75 630 77 678
rect 84 630 86 678
rect 102 630 107 678
rect 114 630 116 678
rect 41 549 44 597
rect 51 549 56 597
rect 246 630 263 678
rect 270 630 280 678
rect 296 630 321 678
rect 328 630 331 678
rect 105 551 107 599
rect 114 551 142 599
rect 158 551 160 599
rect 167 551 177 599
rect 193 551 201 599
rect 208 551 210 599
rect 226 551 263 599
rect 270 551 272 599
rect 386 551 389 599
rect 396 551 406 599
rect 75 425 77 473
rect 84 425 87 473
rect 103 425 107 473
rect 114 425 116 473
rect 136 425 160 473
rect 167 425 175 473
rect 193 425 201 473
rect 208 425 210 473
rect 226 425 263 473
rect 270 425 273 473
rect 350 425 353 473
rect 360 425 366 473
<< ntransistor >>
rect 141 325 148 363
rect 181 325 188 363
rect 222 325 229 363
rect 263 325 270 363
rect 77 255 84 285
rect 141 255 148 285
rect 44 187 51 217
rect 353 255 360 285
rect 141 187 148 217
rect 181 187 188 217
rect 263 187 270 217
rect 321 187 328 217
rect 77 128 84 158
rect 222 128 229 158
rect 263 128 270 158
rect 386 147 393 177
<< ptransistor >>
rect 77 630 84 678
rect 107 630 114 678
rect 44 549 51 597
rect 263 630 270 678
rect 321 630 328 678
rect 107 551 114 599
rect 160 551 167 599
rect 201 551 208 599
rect 263 551 270 599
rect 389 551 396 599
rect 77 425 84 473
rect 107 425 114 473
rect 160 425 167 473
rect 201 425 208 473
rect 263 425 270 473
rect 353 425 360 473
<< polycontact >>
rect 142 682 158 698
rect 192 632 208 648
rect 380 662 396 678
rect 344 526 360 542
rect 316 503 332 519
rect 35 372 51 388
rect 160 399 176 415
rect 263 399 279 415
rect 73 312 89 328
rect 265 229 281 245
rect 344 325 360 363
rect 213 187 229 217
rect 321 147 337 177
rect 370 187 386 217
rect 136 108 152 124
rect 177 108 194 125
<< ndiffcontact >>
rect 120 325 136 363
rect 195 325 211 363
rect 275 325 291 363
rect 56 255 72 285
rect 159 255 175 285
rect 26 187 42 217
rect 56 187 72 217
rect 335 255 351 285
rect 366 255 382 285
rect 123 187 139 217
rect 191 187 207 217
rect 239 187 255 217
rect 332 187 348 217
rect 56 128 72 158
rect 89 128 105 158
rect 204 128 220 158
rect 274 128 290 158
rect 367 147 383 177
rect 396 147 412 177
<< pdiffcontact >>
rect 59 630 75 678
rect 86 630 102 678
rect 116 630 132 678
rect 25 549 41 597
rect 56 549 72 597
rect 230 630 246 678
rect 280 630 296 678
rect 331 630 347 678
rect 89 551 105 599
rect 142 551 158 599
rect 177 551 193 599
rect 210 551 226 599
rect 272 551 288 599
rect 370 551 386 599
rect 406 551 422 599
rect 59 425 75 473
rect 87 425 103 473
rect 116 425 136 473
rect 175 425 193 473
rect 210 425 226 473
rect 273 425 289 473
rect 334 425 350 473
rect 366 425 383 473
<< psubstratetap >>
rect 230 77 247 94
<< nsubstratetap >>
rect 240 714 257 731
<< metal1 >>
rect 0 769 429 779
rect 0 746 319 756
rect 335 746 429 756
rect 0 731 429 733
rect 0 714 240 731
rect 257 714 429 731
rect 0 708 429 714
rect 25 621 41 708
rect 59 678 75 708
rect 86 688 142 698
rect 86 678 102 688
rect 280 688 380 698
rect 280 678 296 688
rect 380 678 396 682
rect 25 620 42 621
rect 116 620 132 630
rect 25 608 132 620
rect 142 632 192 642
rect 25 597 41 608
rect 89 599 105 608
rect 25 498 41 549
rect 142 599 158 632
rect 230 620 246 630
rect 331 620 347 630
rect 406 620 422 708
rect 177 610 422 620
rect 177 599 193 610
rect 272 599 288 610
rect 406 599 422 610
rect 56 536 72 549
rect 142 536 158 551
rect 56 526 158 536
rect 210 541 226 551
rect 210 531 344 541
rect 116 503 290 513
rect 306 503 316 513
rect 370 513 386 551
rect 332 503 386 513
rect 25 488 103 498
rect 87 473 103 488
rect 116 473 136 503
rect 406 493 422 551
rect 175 483 289 493
rect 175 473 193 483
rect 273 473 289 483
rect 334 483 422 493
rect 334 473 350 483
rect 289 425 334 473
rect 59 415 75 425
rect 210 415 226 425
rect 366 415 383 425
rect 59 405 160 415
rect 176 405 226 415
rect 279 405 383 415
rect 14 375 35 385
rect 74 377 211 389
rect 74 350 87 377
rect 195 363 211 377
rect 26 338 87 350
rect 26 285 42 338
rect 73 311 89 312
rect 291 325 344 363
rect 120 315 136 325
rect 120 305 412 315
rect 26 255 56 285
rect 175 275 335 285
rect 26 217 42 255
rect 56 244 72 255
rect 366 245 382 255
rect 56 232 255 244
rect 239 217 255 232
rect 281 229 382 245
rect 72 187 123 217
rect 207 187 213 217
rect 348 187 370 217
rect 26 158 42 187
rect 396 177 412 305
rect 26 128 56 158
rect 105 148 204 158
rect 337 147 367 177
rect 26 98 44 128
rect 135 108 136 124
rect 274 118 290 128
rect 194 108 290 118
rect 14 94 429 98
rect 14 77 230 94
rect 247 77 429 94
rect 14 73 429 77
rect 14 50 73 60
rect 89 50 429 60
rect 14 27 429 37
rect 14 4 119 14
rect 135 4 429 14
<< m2contact >>
rect 319 743 335 759
rect 380 682 396 698
rect 290 503 306 519
rect 73 295 89 311
rect 119 108 135 124
rect 73 47 89 63
rect 119 0 135 16
<< metal2 >>
rect 292 519 304 780
rect 321 759 333 780
rect 321 698 333 743
rect 321 682 380 698
rect 73 63 89 295
rect 119 16 135 108
rect 292 4 304 503
rect 321 4 333 682
<< labels >>
rlabel metal1 14 73 14 98 3 GND!
rlabel metal1 14 4 14 14 3 nRst
rlabel metal1 14 27 14 37 3 Test
rlabel metal1 14 50 14 60 3 Clk
rlabel metal1 0 746 0 756 3 Q
rlabel metal1 0 708 0 733 3 Vdd!
rlabel metal1 0 769 0 779 3 ScanReturn
rlabel metal2 321 4 333 4 1 Q
rlabel metal2 292 4 304 4 1 nQ
rlabel metal1 14 375 14 385 3 D
rlabel metal2 321 780 333 780 5 Q
rlabel metal2 292 780 304 780 5 nQ
<< end >>
