magic
tech c035u
timestamp 1385919140
<< nwell >>
rect 0 403 120 747
<< polysilicon >>
rect 63 532 70 540
rect 33 463 40 471
rect 33 405 40 415
rect 33 353 40 389
rect 63 379 70 484
rect 33 315 40 323
rect 63 310 70 363
rect 63 271 70 280
<< ndiffusion >>
rect 31 323 33 353
rect 40 323 42 353
rect 61 280 63 310
rect 70 309 96 310
rect 70 280 80 309
<< pdiffusion >>
rect 58 484 63 532
rect 70 484 80 532
rect 31 415 33 463
rect 40 415 42 463
<< pohmic >>
rect 0 77 6 87
rect 22 77 34 87
rect 50 77 62 87
rect 78 77 90 87
rect 106 77 120 87
<< nohmic >>
rect 0 737 6 747
rect 23 737 35 747
rect 52 737 64 747
rect 81 737 93 747
rect 110 737 120 747
<< ntransistor >>
rect 33 323 40 353
rect 63 280 70 310
<< ptransistor >>
rect 63 484 70 532
rect 33 415 40 463
<< polycontact >>
rect 32 389 48 405
rect 54 363 70 379
<< ndiffcontact >>
rect 15 323 31 353
rect 42 323 58 353
rect 45 280 61 310
rect 80 280 96 309
<< pdiffcontact >>
rect 42 484 58 532
rect 80 484 96 532
rect 15 415 31 463
rect 42 415 58 463
<< psubstratetap >>
rect 6 77 22 93
rect 34 77 50 93
rect 62 77 78 93
rect 90 77 106 93
<< nsubstratetap >>
rect 6 731 23 747
rect 35 731 52 747
rect 64 731 81 747
rect 93 731 110 747
<< metal1 >>
rect 0 783 120 793
rect 0 760 120 770
rect 0 731 6 747
rect 23 731 35 747
rect 52 731 64 747
rect 81 731 93 747
rect 110 731 120 747
rect 0 722 120 731
rect 42 532 58 722
rect 15 484 42 532
rect 15 463 31 484
rect 31 389 32 405
rect 58 379 68 463
rect 80 405 96 484
rect 58 323 68 363
rect 15 310 31 323
rect 15 280 45 310
rect 45 102 61 280
rect 80 309 96 389
rect 80 279 96 280
rect 0 93 120 102
rect 0 77 6 93
rect 22 77 34 93
rect 50 77 62 93
rect 78 77 90 93
rect 106 77 120 93
rect 0 54 120 64
rect 0 31 120 41
rect 0 8 120 18
<< m2contact >>
rect 15 389 31 405
rect 80 389 96 405
<< metal2 >>
rect 15 405 31 800
rect 15 1 31 389
rect 80 405 96 800
rect 80 1 96 389
<< labels >>
rlabel metal1 0 77 0 102 3 GND!
rlabel metal1 0 54 0 64 3 Clock
rlabel metal1 0 31 0 41 3 Test
rlabel metal1 0 8 0 18 2 nReset
rlabel metal1 120 8 120 18 8 nReset
rlabel metal1 120 31 120 41 7 Test
rlabel metal1 120 54 120 64 7 Clock
rlabel metal1 120 77 120 102 7 GND!
rlabel metal2 15 1 31 1 1 A
rlabel metal2 80 1 96 1 1 Y
rlabel metal1 0 783 0 793 4 ScanReturn
rlabel metal1 0 760 0 770 3 Scan
rlabel metal1 0 722 0 747 3 Vdd!
rlabel metal1 120 722 120 747 7 Vdd!
rlabel metal1 120 760 120 770 7 Scan
rlabel metal1 120 783 120 793 6 ScanReturn
rlabel metal2 15 800 31 800 5 A
rlabel metal2 80 800 96 800 5 Y
<< end >>
