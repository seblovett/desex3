magic
tech c035u
timestamp 1385926013
<< nwell >>
rect 0 402 192 746
<< polysilicon >>
rect 29 691 36 699
rect 59 691 66 699
rect 88 691 95 699
rect 115 691 122 699
rect 146 691 153 699
rect 29 612 36 643
rect 59 599 66 643
rect 29 347 36 564
rect 59 347 66 583
rect 88 573 95 643
rect 115 591 122 643
rect 146 633 153 643
rect 149 617 153 633
rect 115 575 116 591
rect 88 347 95 557
rect 115 347 122 575
rect 146 393 153 617
rect 148 377 153 393
rect 29 282 36 317
rect 59 278 66 317
rect 88 309 95 317
rect 115 309 122 317
rect 146 282 153 377
rect 29 242 36 252
rect 146 244 153 252
rect 29 226 37 242
<< ndiffusion >>
rect 27 317 29 347
rect 36 317 38 347
rect 54 317 59 347
rect 66 317 88 347
rect 95 317 97 347
rect 113 317 115 347
rect 122 317 124 347
rect 27 252 29 282
rect 36 252 38 282
rect 144 252 146 282
rect 153 252 155 282
<< pdiffusion >>
rect 27 643 29 691
rect 36 643 38 691
rect 54 643 59 691
rect 66 643 68 691
rect 84 643 88 691
rect 95 643 97 691
rect 113 643 115 691
rect 122 643 125 691
rect 141 643 146 691
rect 153 643 156 691
rect 27 564 29 612
rect 36 564 38 612
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 192 86
rect 0 76 192 79
<< nohmic >>
rect 0 743 192 746
rect 0 736 8 743
rect 24 736 36 743
rect 52 736 64 743
rect 80 736 92 743
rect 108 736 120 743
rect 136 736 148 743
rect 164 736 192 743
<< ntransistor >>
rect 29 317 36 347
rect 59 317 66 347
rect 88 317 95 347
rect 115 317 122 347
rect 29 252 36 282
rect 146 252 153 282
<< ptransistor >>
rect 29 643 36 691
rect 59 643 66 691
rect 88 643 95 691
rect 115 643 122 691
rect 146 643 153 691
rect 29 564 36 612
<< polycontact >>
rect 59 583 75 599
rect 133 617 149 633
rect 116 575 132 591
rect 84 557 100 573
rect 132 377 148 393
rect 59 262 75 278
rect 37 226 53 242
<< ndiffcontact >>
rect 11 317 27 347
rect 38 317 54 347
rect 97 317 113 347
rect 124 317 140 347
rect 11 252 27 282
rect 38 252 54 282
rect 128 252 144 282
rect 155 252 175 282
<< pdiffcontact >>
rect 11 643 27 691
rect 38 643 54 691
rect 68 643 84 691
rect 97 643 113 691
rect 125 643 141 691
rect 156 643 176 691
rect 11 564 27 612
rect 38 564 54 612
<< psubstratetap >>
rect 6 79 22 95
rect 34 79 50 95
rect 62 79 78 95
rect 90 79 106 95
rect 118 79 134 95
rect 146 79 162 95
<< nsubstratetap >>
rect 8 727 24 743
rect 36 727 52 743
rect 64 727 80 743
rect 92 727 108 743
rect 120 727 136 743
rect 148 727 164 743
<< metal1 >>
rect 0 782 192 792
rect 0 759 118 769
rect 0 743 192 746
rect 0 727 8 743
rect 24 727 36 743
rect 52 727 64 743
rect 80 727 92 743
rect 108 727 120 743
rect 136 727 148 743
rect 164 727 192 743
rect 0 721 192 727
rect 11 691 27 721
rect 41 701 110 711
rect 41 691 51 701
rect 100 691 110 701
rect 125 691 141 721
rect 11 612 27 643
rect 71 629 81 643
rect 71 619 133 629
rect 54 583 59 599
rect 41 380 132 390
rect 41 347 51 380
rect 159 385 169 643
rect 159 375 192 385
rect 73 357 137 367
rect 14 307 24 317
rect 73 307 83 357
rect 127 347 137 357
rect 14 297 83 307
rect 54 262 59 278
rect 11 101 27 252
rect 97 101 113 317
rect 159 282 169 375
rect 128 101 144 252
rect 0 95 192 101
rect 0 79 6 95
rect 22 79 34 95
rect 50 79 62 95
rect 78 79 90 95
rect 106 79 118 95
rect 134 79 146 95
rect 162 79 192 95
rect 0 76 192 79
rect 0 53 192 63
rect 0 30 39 40
rect 53 30 192 40
rect 0 7 192 17
<< m2contact >>
rect 118 757 132 771
rect 118 591 132 605
rect 85 543 99 557
rect 39 212 53 226
rect 39 28 53 42
<< metal2 >>
rect 96 557 108 799
rect 119 605 131 757
rect 99 543 108 557
rect 40 42 52 212
rect 96 0 108 543
<< labels >>
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal2 96 799 108 799 5 D
rlabel metal1 0 76 0 101 1 GND!
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 3 Clock
rlabel metal2 96 0 108 0 1 D
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 192 782 192 792 6 ScanReturn
rlabel metal1 192 53 192 63 7 Clock
rlabel metal1 192 30 192 40 7 Test
rlabel metal1 192 7 192 17 8 nReset
rlabel metal1 192 76 192 101 7 GND!
rlabel metal1 192 721 192 746 7 Vdd!
rlabel metal1 192 375 192 385 7 M
<< end >>
