magic
tech c035u
timestamp 1386541191
<< metal1 >>
rect 1951 840 1971 850
rect 0 802 31 827
rect 0 157 31 182
rect 1951 134 1963 144
rect 1951 111 2019 121
rect 1951 88 1986 98
rect 1556 65 1986 75
rect 1796 43 1962 53
rect 1676 17 2019 27
<< m2contact >>
rect 1971 837 1985 851
rect 1963 131 1977 145
rect 2019 109 2033 123
rect 1986 87 2000 101
rect 1542 63 1556 77
rect 1986 63 2000 77
rect 1782 41 1796 55
rect 1962 41 1976 55
rect 1662 15 1676 29
rect 2019 15 2033 29
<< metal2 >>
rect 55 956 1435 968
rect 55 880 67 956
rect 103 934 1315 946
rect 103 880 115 934
rect 583 912 1147 924
rect 583 880 595 912
rect 631 890 907 902
rect 631 880 643 890
rect 775 880 787 890
rect 895 880 907 890
rect 1015 880 1027 912
rect 1135 880 1147 912
rect 1303 880 1315 934
rect 1423 880 1435 956
rect 1903 894 1984 906
rect 1903 880 1915 894
rect 1972 851 1984 894
rect 55 0 67 81
rect 103 0 115 81
rect 583 0 595 81
rect 631 0 643 81
rect 1255 0 1267 81
rect 1375 0 1387 81
rect 1495 0 1507 81
rect 1543 77 1555 81
rect 1543 0 1555 63
rect 1615 0 1627 81
rect 1663 29 1675 81
rect 1663 0 1675 15
rect 1735 0 1747 81
rect 1783 55 1795 81
rect 1783 0 1795 41
rect 1855 0 1867 81
rect 1964 55 1976 131
rect 1987 77 1999 87
rect 2020 29 2032 109
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 31 0 1 81
box 0 0 720 799
use inv inv_0
timestamp 1386238110
transform 1 0 751 0 1 81
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 871 0 1 81
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 991 0 1 81
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 1111 0 1 81
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 1231 0 1 81
box 0 0 120 799
use inv inv_5
timestamp 1386238110
transform 1 0 1351 0 1 81
box 0 0 120 799
use inv inv_6
timestamp 1386238110
transform 1 0 1471 0 1 81
box 0 0 120 799
use inv inv_7
timestamp 1386238110
transform 1 0 1591 0 1 81
box 0 0 120 799
use inv inv_8
timestamp 1386238110
transform 1 0 1711 0 1 81
box 0 0 120 799
use inv inv_9
timestamp 1386238110
transform 1 0 1831 0 1 81
box 0 0 120 799
<< labels >>
rlabel metal2 1735 0 1747 0 1 nClock
rlabel metal2 1855 0 1867 0 1 nSDI
rlabel metal2 1375 0 1387 0 1 nD
rlabel metal2 1255 0 1267 0 1 nLoad
rlabel metal2 103 0 115 0 1 Load
rlabel metal2 55 0 67 0 1 D
rlabel metal2 631 0 643 0 1 Q
rlabel metal2 583 0 595 0 1 nQ
rlabel metal2 1663 0 1675 0 1 Test
rlabel metal2 1783 0 1795 0 1 Clock
rlabel metal1 0 157 0 182 3 GND!
rlabel metal1 0 802 0 827 3 Vdd!
rlabel metal2 1615 0 1627 0 1 nTest
rlabel metal2 1543 0 1555 0 1 nReset
rlabel metal2 1495 0 1507 0 1 nnReset
<< end >>
