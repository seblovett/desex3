magic
tech c035u
timestamp 1385058125
<< error_p >>
rect 352 488 357 490
rect 1336 86 1337 92
<< nwell >>
rect 202 524 1442 736
rect 202 522 1332 524
rect 202 491 1331 522
rect 202 490 1318 491
rect 202 488 329 490
rect 352 398 644 490
rect 689 398 981 490
rect 1026 398 1318 490
rect 405 397 451 398
rect 742 397 788 398
rect 1079 397 1125 398
<< polysilicon >>
rect 538 688 545 696
rect 565 688 572 696
rect 592 688 599 696
rect 619 688 626 696
rect 875 688 882 696
rect 902 688 909 696
rect 929 688 936 696
rect 956 688 963 696
rect 1212 688 1219 696
rect 1239 688 1246 696
rect 1266 688 1273 696
rect 1293 688 1300 696
rect 480 610 487 618
rect 507 610 514 618
rect 370 456 377 584
rect 425 555 432 563
rect 817 610 824 618
rect 844 610 851 618
rect 707 456 714 584
rect 762 555 769 563
rect 1154 610 1161 618
rect 1181 610 1188 618
rect 1044 456 1051 584
rect 1099 555 1106 563
rect 1394 637 1396 653
rect 1389 592 1396 637
rect 1389 496 1396 544
rect 1389 458 1396 466
rect 370 384 377 398
rect 425 384 432 398
rect 480 385 487 398
rect 375 368 377 384
rect 430 368 432 384
rect 485 381 487 385
rect 507 381 514 398
rect 538 385 545 398
rect 485 374 514 381
rect 485 369 487 374
rect 543 381 545 385
rect 565 381 572 398
rect 592 381 599 398
rect 619 381 626 398
rect 707 384 714 398
rect 762 384 769 398
rect 817 385 824 398
rect 543 374 626 381
rect 543 369 545 374
rect 370 358 377 368
rect 425 358 432 368
rect 480 358 487 369
rect 538 358 545 369
rect 565 358 572 374
rect 712 368 714 384
rect 767 368 769 384
rect 822 381 824 385
rect 844 381 851 398
rect 875 385 882 398
rect 822 374 851 381
rect 822 369 824 374
rect 880 381 882 385
rect 902 381 909 398
rect 929 381 936 398
rect 956 381 963 398
rect 1044 384 1051 398
rect 1099 384 1106 398
rect 1154 385 1161 398
rect 880 374 963 381
rect 880 369 882 374
rect 707 358 714 368
rect 762 358 769 368
rect 817 358 824 369
rect 875 358 882 369
rect 902 358 909 374
rect 1049 368 1051 384
rect 1104 368 1106 384
rect 1159 381 1161 385
rect 1181 381 1188 398
rect 1212 385 1219 398
rect 1159 374 1188 381
rect 1159 369 1161 374
rect 1217 381 1219 385
rect 1239 381 1246 398
rect 1266 381 1273 398
rect 1293 381 1300 398
rect 1217 374 1300 381
rect 1217 369 1219 374
rect 1044 358 1051 368
rect 1099 358 1106 368
rect 1154 358 1161 369
rect 1212 358 1219 369
rect 1239 358 1246 374
rect 370 330 377 338
rect 425 296 432 304
rect 480 204 487 212
rect 707 330 714 338
rect 762 296 769 304
rect 817 204 824 212
rect 1044 330 1051 338
rect 1099 296 1106 304
rect 1154 204 1161 212
rect 538 150 545 158
rect 565 150 572 158
rect 875 150 882 158
rect 902 150 909 158
rect 1212 150 1219 158
rect 1239 150 1246 158
<< ndiffusion >>
rect 1387 466 1389 496
rect 1396 466 1398 496
rect 368 338 370 358
rect 377 338 379 358
rect 423 304 425 358
rect 432 304 434 358
rect 478 212 480 358
rect 487 212 489 358
rect 536 158 538 358
rect 545 158 547 358
rect 563 158 565 358
rect 572 158 574 358
rect 705 338 707 358
rect 714 338 716 358
rect 760 304 762 358
rect 769 304 771 358
rect 815 212 817 358
rect 824 212 826 358
rect 873 158 875 358
rect 882 158 884 358
rect 900 158 902 358
rect 909 158 911 358
rect 1042 338 1044 358
rect 1051 338 1053 358
rect 1097 304 1099 358
rect 1106 304 1108 358
rect 1152 212 1154 358
rect 1161 212 1163 358
rect 1210 158 1212 358
rect 1219 158 1221 358
rect 1237 158 1239 358
rect 1246 158 1248 358
<< pdiffusion >>
rect 368 398 370 456
rect 377 398 379 456
rect 423 398 425 555
rect 432 398 434 555
rect 478 398 480 610
rect 487 398 489 610
rect 505 398 507 610
rect 514 398 516 610
rect 536 398 538 688
rect 545 398 547 688
rect 563 398 565 688
rect 572 398 574 688
rect 590 398 592 688
rect 599 398 601 688
rect 617 398 619 688
rect 626 398 628 688
rect 705 398 707 456
rect 714 398 716 456
rect 760 398 762 555
rect 769 398 771 555
rect 815 398 817 610
rect 824 398 826 610
rect 842 398 844 610
rect 851 398 853 610
rect 873 398 875 688
rect 882 398 884 688
rect 900 398 902 688
rect 909 398 911 688
rect 927 398 929 688
rect 936 398 938 688
rect 954 398 956 688
rect 963 398 965 688
rect 1042 398 1044 456
rect 1051 398 1053 456
rect 1097 398 1099 555
rect 1106 398 1108 555
rect 1152 398 1154 610
rect 1161 398 1163 610
rect 1179 398 1181 610
rect 1188 398 1190 610
rect 1210 398 1212 688
rect 1219 398 1221 688
rect 1237 398 1239 688
rect 1246 398 1248 688
rect 1264 398 1266 688
rect 1273 398 1275 688
rect 1291 398 1293 688
rect 1300 398 1302 688
rect 1387 544 1389 592
rect 1396 544 1398 592
<< pohmic >>
rect 320 76 326 86
rect 342 76 354 86
rect 370 76 382 86
rect 398 76 410 86
rect 426 76 438 86
rect 454 76 466 86
rect 482 76 494 86
rect 510 76 522 86
rect 538 76 550 86
rect 567 76 579 86
rect 595 76 607 86
rect 623 76 635 86
rect 651 76 663 86
rect 679 76 691 86
rect 707 76 719 86
rect 735 76 747 86
rect 763 76 775 86
rect 791 76 803 86
rect 819 76 831 86
rect 847 76 859 86
rect 875 76 887 86
rect 904 76 916 86
rect 932 76 944 86
rect 960 76 972 86
rect 988 76 1000 86
rect 1016 76 1028 86
rect 1044 76 1056 86
rect 1072 76 1084 86
rect 1100 76 1112 86
rect 1128 76 1140 86
rect 1156 76 1168 86
rect 1184 76 1196 86
rect 1212 76 1224 86
rect 1241 76 1253 86
rect 1269 76 1281 86
rect 1297 76 1309 86
rect 1325 76 1336 86
rect 1352 76 1364 86
rect 1380 76 1392 86
rect 1408 76 1420 86
rect 1436 76 1442 86
<< nohmic >>
rect 202 726 214 736
rect 230 726 242 736
rect 258 726 270 736
rect 286 726 298 736
rect 314 726 326 736
rect 342 726 354 736
rect 370 726 382 736
rect 398 726 410 736
rect 426 726 438 736
rect 454 726 466 736
rect 482 726 494 736
rect 510 726 522 736
rect 538 726 550 736
rect 567 726 579 736
rect 595 726 607 736
rect 623 726 635 736
rect 651 726 663 736
rect 679 726 691 736
rect 707 726 719 736
rect 735 726 747 736
rect 763 726 775 736
rect 791 726 803 736
rect 819 726 831 736
rect 847 726 859 736
rect 875 726 887 736
rect 904 726 916 736
rect 932 726 944 736
rect 960 726 972 736
rect 988 726 1000 736
rect 1016 726 1028 736
rect 1044 726 1056 736
rect 1072 726 1084 736
rect 1100 726 1112 736
rect 1128 726 1140 736
rect 1156 726 1168 736
rect 1184 726 1196 736
rect 1212 726 1224 736
rect 1241 726 1253 736
rect 1269 726 1281 736
rect 1297 726 1309 736
rect 1325 726 1337 736
rect 1353 726 1365 736
rect 1381 726 1393 736
rect 1409 726 1421 736
rect 1437 726 1442 736
<< ntransistor >>
rect 1389 466 1396 496
rect 370 338 377 358
rect 425 304 432 358
rect 480 212 487 358
rect 538 158 545 358
rect 565 158 572 358
rect 707 338 714 358
rect 762 304 769 358
rect 817 212 824 358
rect 875 158 882 358
rect 902 158 909 358
rect 1044 338 1051 358
rect 1099 304 1106 358
rect 1154 212 1161 358
rect 1212 158 1219 358
rect 1239 158 1246 358
<< ptransistor >>
rect 370 398 377 456
rect 425 398 432 555
rect 480 398 487 610
rect 507 398 514 610
rect 538 398 545 688
rect 565 398 572 688
rect 592 398 599 688
rect 619 398 626 688
rect 707 398 714 456
rect 762 398 769 555
rect 817 398 824 610
rect 844 398 851 610
rect 875 398 882 688
rect 902 398 909 688
rect 929 398 936 688
rect 956 398 963 688
rect 1044 398 1051 456
rect 1099 398 1106 555
rect 1154 398 1161 610
rect 1181 398 1188 610
rect 1212 398 1219 688
rect 1239 398 1246 688
rect 1266 398 1273 688
rect 1293 398 1300 688
rect 1389 544 1396 592
<< polycontact >>
rect 1378 637 1394 653
rect 359 368 375 384
rect 414 368 430 384
rect 469 369 485 385
rect 527 369 543 385
rect 696 368 712 384
rect 751 368 767 384
rect 806 369 822 385
rect 864 369 880 385
rect 1033 368 1049 384
rect 1088 368 1104 384
rect 1143 369 1159 385
rect 1201 369 1217 385
<< ndiffcontact >>
rect 1371 466 1387 496
rect 1398 466 1414 496
rect 352 338 368 358
rect 379 338 395 358
rect 407 304 423 358
rect 434 304 450 358
rect 462 212 478 358
rect 489 212 505 358
rect 520 158 536 358
rect 547 158 563 358
rect 574 158 590 358
rect 689 338 705 358
rect 716 338 732 358
rect 744 304 760 358
rect 771 304 787 358
rect 799 212 815 358
rect 826 212 842 358
rect 857 158 873 358
rect 884 158 900 358
rect 911 158 927 358
rect 1026 338 1042 358
rect 1053 338 1069 358
rect 1081 304 1097 358
rect 1108 304 1124 358
rect 1136 212 1152 358
rect 1163 212 1179 358
rect 1194 158 1210 358
rect 1221 158 1237 358
rect 1248 158 1264 358
<< pdiffcontact >>
rect 519 610 536 688
rect 352 398 368 456
rect 379 398 395 456
rect 407 398 423 555
rect 434 398 450 555
rect 462 398 478 610
rect 489 398 505 610
rect 516 398 536 610
rect 547 398 563 688
rect 574 398 590 688
rect 601 398 617 688
rect 628 398 644 688
rect 856 610 873 688
rect 689 398 705 456
rect 716 398 732 456
rect 744 398 760 555
rect 771 398 787 555
rect 799 398 815 610
rect 826 398 842 610
rect 853 398 873 610
rect 884 398 900 688
rect 911 398 927 688
rect 938 398 954 688
rect 965 398 981 688
rect 1193 610 1210 688
rect 1026 398 1042 456
rect 1053 398 1069 456
rect 1081 398 1097 555
rect 1108 398 1124 555
rect 1136 398 1152 610
rect 1163 398 1179 610
rect 1190 398 1210 610
rect 1221 398 1237 688
rect 1248 398 1264 688
rect 1275 398 1291 688
rect 1302 398 1318 688
rect 1371 544 1387 592
rect 1398 544 1414 592
<< psubstratetap >>
rect 326 76 342 92
rect 354 76 370 92
rect 382 76 398 92
rect 410 76 426 92
rect 438 76 454 92
rect 466 76 482 92
rect 494 76 510 92
rect 522 76 538 92
rect 550 76 567 92
rect 579 76 595 92
rect 607 76 623 92
rect 635 76 651 92
rect 663 76 679 92
rect 691 76 707 92
rect 719 76 735 92
rect 747 76 763 92
rect 775 76 791 92
rect 803 76 819 92
rect 831 76 847 92
rect 859 76 875 92
rect 887 76 904 92
rect 916 76 932 92
rect 944 76 960 92
rect 972 76 988 92
rect 1000 76 1016 92
rect 1028 76 1044 92
rect 1056 76 1072 92
rect 1084 76 1100 92
rect 1112 76 1128 92
rect 1140 76 1156 92
rect 1168 76 1184 92
rect 1196 76 1212 92
rect 1224 76 1241 92
rect 1253 76 1269 92
rect 1281 76 1297 92
rect 1309 76 1325 92
rect 1336 76 1352 92
rect 1364 76 1380 92
rect 1392 76 1408 92
rect 1420 76 1436 92
<< nsubstratetap >>
rect 214 720 230 736
rect 242 720 258 736
rect 270 720 286 736
rect 298 720 314 736
rect 326 720 342 736
rect 354 720 370 736
rect 382 720 398 736
rect 410 720 426 736
rect 438 720 454 736
rect 466 720 482 736
rect 494 720 510 736
rect 522 720 538 736
rect 550 720 567 736
rect 579 720 595 736
rect 607 720 623 736
rect 635 720 651 736
rect 663 720 679 736
rect 691 720 707 736
rect 719 720 735 736
rect 747 720 763 736
rect 775 720 791 736
rect 803 720 819 736
rect 831 720 847 736
rect 859 720 875 736
rect 887 720 904 736
rect 916 720 932 736
rect 944 720 960 736
rect 972 720 988 736
rect 1000 720 1016 736
rect 1028 720 1044 736
rect 1056 720 1072 736
rect 1084 720 1100 736
rect 1112 720 1128 736
rect 1140 720 1156 736
rect 1168 720 1184 736
rect 1196 720 1212 736
rect 1224 720 1241 736
rect 1253 720 1269 736
rect 1281 720 1297 736
rect 1309 720 1325 736
rect 1337 720 1353 736
rect 1365 720 1381 736
rect 1393 720 1409 736
rect 1421 720 1437 736
<< metal1 >>
rect 236 772 1356 782
rect 1400 772 1442 782
rect 236 749 1442 759
rect 200 720 214 736
rect 230 720 242 736
rect 258 720 270 736
rect 286 720 298 736
rect 314 720 326 736
rect 342 720 354 736
rect 370 720 382 736
rect 398 720 410 736
rect 426 720 438 736
rect 454 720 466 736
rect 482 720 494 736
rect 510 720 522 736
rect 538 720 550 736
rect 567 720 579 736
rect 595 720 607 736
rect 623 720 635 736
rect 651 720 663 736
rect 679 720 691 736
rect 707 720 719 736
rect 735 720 747 736
rect 763 720 775 736
rect 791 720 803 736
rect 819 720 831 736
rect 847 720 859 736
rect 875 720 887 736
rect 904 720 916 736
rect 932 720 944 736
rect 960 720 972 736
rect 988 720 1000 736
rect 1016 720 1028 736
rect 1044 720 1056 736
rect 1072 720 1084 736
rect 1100 720 1112 736
rect 1128 720 1140 736
rect 1156 720 1168 736
rect 1184 720 1196 736
rect 1212 720 1224 736
rect 1241 720 1253 736
rect 1269 720 1281 736
rect 1297 720 1309 736
rect 1325 720 1337 736
rect 1353 720 1365 736
rect 1381 720 1393 736
rect 1409 720 1421 736
rect 1437 720 1442 736
rect 200 711 1442 720
rect 352 456 368 711
rect 407 555 423 711
rect 462 610 478 711
rect 516 688 536 711
rect 574 688 590 711
rect 628 688 644 711
rect 516 610 519 688
rect 689 456 705 711
rect 744 555 760 711
rect 799 610 815 711
rect 853 688 873 711
rect 911 688 927 711
rect 965 688 981 711
rect 853 610 856 688
rect 1026 456 1042 711
rect 1081 555 1097 711
rect 1136 610 1152 711
rect 1190 688 1210 711
rect 1248 688 1264 711
rect 1302 688 1318 711
rect 1190 610 1193 688
rect 1380 653 1394 659
rect 1404 592 1414 711
rect 1371 496 1381 544
rect 284 371 359 381
rect 385 381 395 398
rect 385 371 414 381
rect 385 358 395 371
rect 440 382 450 398
rect 440 372 469 382
rect 440 358 450 372
rect 495 382 505 398
rect 495 372 527 382
rect 495 358 505 372
rect 553 383 563 398
rect 607 385 617 398
rect 553 373 606 383
rect 553 358 563 373
rect 667 371 696 381
rect 722 381 732 398
rect 722 371 751 381
rect 722 358 732 371
rect 777 382 787 398
rect 777 372 806 382
rect 777 358 787 372
rect 832 382 842 398
rect 832 372 864 382
rect 832 358 842 372
rect 890 383 900 398
rect 944 385 954 398
rect 890 373 944 383
rect 890 358 900 373
rect 1022 371 1033 381
rect 1059 381 1069 398
rect 1059 371 1088 381
rect 1059 358 1069 371
rect 1114 382 1124 398
rect 1114 372 1143 382
rect 1114 358 1124 372
rect 1169 382 1179 398
rect 1169 372 1201 382
rect 1169 358 1179 372
rect 1227 383 1237 398
rect 1281 385 1291 398
rect 1227 373 1279 383
rect 1227 358 1237 373
rect 352 101 368 338
rect 407 101 423 304
rect 462 101 478 212
rect 689 101 705 338
rect 744 101 760 304
rect 799 101 815 212
rect 1026 101 1042 338
rect 1081 101 1097 304
rect 1136 101 1152 212
rect 1398 101 1408 466
rect 320 92 1442 101
rect 320 76 326 92
rect 342 76 354 92
rect 370 76 382 92
rect 398 76 410 92
rect 426 76 438 92
rect 454 76 466 92
rect 482 76 494 92
rect 510 76 522 92
rect 538 76 550 92
rect 567 76 579 92
rect 595 76 607 92
rect 623 76 635 92
rect 651 76 663 92
rect 679 76 691 92
rect 707 76 719 92
rect 735 76 747 92
rect 763 76 775 92
rect 791 76 803 92
rect 819 76 831 92
rect 847 76 859 92
rect 875 76 887 92
rect 904 76 916 92
rect 932 76 944 92
rect 960 76 972 92
rect 988 76 1000 92
rect 1016 76 1028 92
rect 1044 76 1056 92
rect 1072 76 1084 92
rect 1100 76 1112 92
rect 1128 76 1140 92
rect 1156 76 1168 92
rect 1184 76 1196 92
rect 1212 76 1224 92
rect 1241 76 1253 92
rect 1269 76 1281 92
rect 1297 76 1309 92
rect 1325 76 1336 92
rect 1352 76 1364 92
rect 1380 76 1392 92
rect 1408 76 1420 92
rect 1436 76 1442 92
rect 620 53 1442 63
rect 260 30 653 40
rect 959 30 1442 40
rect 308 7 1009 17
rect 1294 7 1442 17
<< m2contact >>
rect 222 771 236 785
rect 1356 771 1370 785
rect 1386 771 1400 785
rect 222 747 236 761
rect 0 711 200 736
rect 1380 659 1394 673
rect 1357 578 1371 592
rect 270 369 284 383
rect 606 371 620 385
rect 653 369 667 383
rect 944 371 958 385
rect 1008 369 1022 383
rect 1279 371 1293 385
rect 606 51 620 65
rect 246 27 260 41
rect 653 28 667 42
rect 945 29 959 43
rect 294 3 308 17
rect 1009 5 1023 19
rect 1280 5 1294 19
<< metal2 >>
rect 0 736 200 790
rect 223 785 235 790
rect 0 -2 200 711
rect 223 -2 235 747
rect 247 41 259 790
rect 271 383 283 790
rect 247 -2 259 27
rect 271 -2 283 369
rect 295 17 307 790
rect 1358 592 1370 771
rect 1386 673 1398 771
rect 1394 659 1398 673
rect 607 65 619 371
rect 654 42 666 369
rect 946 43 958 371
rect 1010 19 1022 369
rect 1281 19 1293 371
rect 295 -2 307 3
<< labels >>
rlabel metal1 1442 711 1442 736 7 Vdd!
rlabel metal1 1442 749 1442 759 7 SDI
rlabel metal1 1442 772 1442 782 7 nSDO
rlabel metal2 0 790 200 790 5 Vdd!
rlabel metal2 223 790 235 790 5 SDO
rlabel metal2 247 790 259 790 5 Test
rlabel metal2 271 790 283 790 5 Clock
rlabel metal2 295 790 307 790 5 nReset
rlabel metal2 247 -2 259 -2 1 Test
rlabel metal2 271 -2 283 -2 1 Clock
rlabel metal2 0 -2 200 -2 1 Vdd!
rlabel metal2 295 -2 307 -2 1 nReset
rlabel metal2 223 -2 235 -2 1 SDI
rlabel metal1 1442 53 1442 63 7 ClockOut
rlabel metal1 1442 30 1442 40 7 TestOut
rlabel metal1 1442 7 1442 17 7 nResetOut
rlabel metal1 1442 76 1442 101 7 GND!
<< end >>
