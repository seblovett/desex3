magic
tech c035u
timestamp 1384456332
<< nwell >>
rect -1 246 465 323
rect 1 220 465 246
rect 2 139 465 220
<< polysilicon >>
rect 87 305 94 313
rect 32 206 39 214
rect 142 289 149 297
rect 169 289 176 297
rect 196 289 203 297
rect 251 293 258 301
rect 278 293 285 301
rect 305 293 312 301
rect 332 293 339 301
rect 359 293 366 301
rect 386 293 393 301
rect 413 293 420 301
rect 440 293 447 301
rect 32 134 39 148
rect 87 134 94 148
rect 142 134 149 148
rect 37 118 39 134
rect 92 118 94 134
rect 147 129 149 134
rect 169 129 176 148
rect 196 129 203 148
rect 251 134 258 148
rect 147 122 203 129
rect 147 118 149 122
rect 32 108 39 118
rect 87 108 94 118
rect 142 108 149 118
rect 169 108 176 122
rect 256 129 258 134
rect 278 129 285 148
rect 305 129 312 148
rect 332 129 339 148
rect 359 129 366 148
rect 386 129 393 148
rect 413 129 420 148
rect 440 131 447 148
rect 438 129 447 131
rect 256 122 447 129
rect 256 118 258 122
rect 251 108 258 118
rect 278 108 285 122
rect 305 108 312 122
rect 332 108 339 122
rect 359 108 366 122
rect 386 108 393 122
rect 413 108 420 122
rect 440 108 447 122
rect 32 80 39 88
rect 87 46 94 54
rect 251 50 258 58
rect 278 50 285 58
rect 305 50 312 58
rect 332 50 339 58
rect 359 50 366 58
rect 386 50 393 58
rect 413 50 420 58
rect 440 50 447 58
rect 142 27 149 35
rect 169 27 176 35
<< ndiffusion >>
rect 30 88 32 108
rect 39 88 41 108
rect 85 54 87 108
rect 94 54 96 108
rect 140 35 142 108
rect 149 35 151 108
rect 167 35 169 108
rect 176 35 178 108
rect 249 58 251 108
rect 258 58 260 108
rect 276 58 278 108
rect 285 58 287 108
rect 303 58 305 108
rect 312 58 314 108
rect 330 58 332 108
rect 339 58 341 108
rect 357 58 359 108
rect 366 58 368 108
rect 384 58 386 108
rect 393 58 395 108
rect 411 58 413 108
rect 420 58 422 108
rect 438 58 440 108
rect 447 58 449 108
<< pdiffusion >>
rect 30 148 32 206
rect 39 148 41 206
rect 85 148 87 305
rect 94 148 96 305
rect 140 148 142 289
rect 149 148 151 289
rect 167 148 169 289
rect 176 148 178 289
rect 194 148 196 289
rect 203 148 205 289
rect 249 148 251 293
rect 258 148 260 293
rect 276 148 278 293
rect 285 148 287 293
rect 303 148 305 293
rect 312 148 314 293
rect 330 148 332 293
rect 339 148 341 293
rect 357 148 359 293
rect 366 148 368 293
rect 384 148 386 293
rect 393 148 395 293
rect 411 148 413 293
rect 420 148 422 293
rect 438 148 440 293
rect 447 148 449 293
<< ntransistor >>
rect 32 88 39 108
rect 87 54 94 108
rect 142 35 149 108
rect 169 35 176 108
rect 251 58 258 108
rect 278 58 285 108
rect 305 58 312 108
rect 332 58 339 108
rect 359 58 366 108
rect 386 58 393 108
rect 413 58 420 108
rect 440 58 447 108
<< ptransistor >>
rect 32 148 39 206
rect 87 148 94 305
rect 142 148 149 289
rect 169 148 176 289
rect 196 148 203 289
rect 251 148 258 293
rect 278 148 285 293
rect 305 148 312 293
rect 332 148 339 293
rect 359 148 366 293
rect 386 148 393 293
rect 413 148 420 293
rect 440 148 447 293
<< polycontact >>
rect 21 118 37 134
rect 76 118 92 134
rect 131 118 147 134
rect 240 118 256 134
<< ndiffcontact >>
rect 14 88 30 108
rect 41 88 57 108
rect 69 54 85 108
rect 96 54 112 108
rect 124 35 140 108
rect 151 35 167 108
rect 178 35 194 108
rect 233 58 249 108
rect 260 58 276 108
rect 287 58 303 108
rect 314 58 330 108
rect 341 58 357 108
rect 368 58 384 108
rect 395 58 411 108
rect 422 58 438 108
rect 449 58 465 108
<< pdiffcontact >>
rect 14 148 30 206
rect 41 148 57 206
rect 69 148 85 305
rect 96 148 112 305
rect 124 148 140 289
rect 151 148 167 289
rect 178 148 194 289
rect 205 148 221 289
rect 233 148 249 293
rect 260 148 276 293
rect 287 148 303 293
rect 314 148 330 293
rect 341 148 357 293
rect 368 148 384 293
rect 395 148 411 293
rect 422 148 438 293
rect 449 148 465 293
<< metal1 >>
rect 0 315 466 340
rect 14 206 30 315
rect 69 305 85 315
rect 124 289 140 315
rect 178 289 194 315
rect 233 293 249 315
rect 287 293 303 315
rect 341 293 357 315
rect 395 293 411 315
rect 449 293 465 315
rect -1 119 21 129
rect 47 131 57 148
rect 47 121 76 131
rect 47 108 57 121
rect 102 131 112 148
rect 102 121 131 131
rect 102 108 112 121
rect 157 131 167 148
rect 211 131 221 148
rect 157 121 240 131
rect 157 108 167 121
rect 266 131 276 148
rect 320 131 330 148
rect 374 131 384 148
rect 428 131 438 148
rect 266 121 459 131
rect 266 108 276 121
rect 320 108 330 121
rect 374 108 384 121
rect 428 108 438 121
rect 14 25 30 88
rect 69 25 85 54
rect 124 25 140 35
rect 178 25 194 35
rect 233 25 249 58
rect 287 25 303 58
rect 341 25 357 58
rect 395 25 411 58
rect 449 25 465 58
rect -1 0 466 25
<< labels >>
rlabel metal1 466 315 466 340 7 Vdd!
rlabel metal1 466 0 466 25 7 GND!
<< end >>
