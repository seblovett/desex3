magic
tech c035u
timestamp 1385636469
<< nwell >>
rect 0 402 603 746
<< polysilicon >>
rect 29 691 36 699
rect 59 691 66 699
rect 88 691 95 699
rect 115 691 122 699
rect 146 691 153 699
rect 251 691 258 719
rect 281 691 288 719
rect 332 704 399 711
rect 29 612 36 643
rect 59 599 66 643
rect 29 347 36 564
rect 59 347 66 583
rect 88 573 95 643
rect 115 591 122 643
rect 146 633 153 643
rect 149 617 153 633
rect 115 575 116 591
rect 88 347 95 557
rect 115 347 122 575
rect 146 393 153 617
rect 218 610 225 621
rect 148 377 153 393
rect 218 388 225 562
rect 251 486 258 643
rect 281 612 288 643
rect 334 612 341 623
rect 375 612 382 645
rect 392 624 399 704
rect 437 691 444 719
rect 495 691 502 719
rect 437 624 444 643
rect 392 617 444 624
rect 437 612 444 617
rect 281 486 288 564
rect 334 486 341 564
rect 375 486 382 564
rect 437 486 444 564
rect 495 532 502 643
rect 563 612 570 675
rect 29 282 36 317
rect 59 278 66 317
rect 88 309 95 317
rect 115 309 122 317
rect 146 282 153 377
rect 29 242 36 252
rect 146 244 153 252
rect 29 226 37 242
rect 218 220 225 372
rect 251 331 258 438
rect 281 402 288 438
rect 334 428 341 438
rect 350 412 362 419
rect 281 395 322 402
rect 315 366 322 395
rect 355 366 362 412
rect 375 410 382 438
rect 437 428 444 438
rect 375 403 403 410
rect 396 366 403 403
rect 437 366 444 412
rect 251 288 258 315
rect 315 288 322 328
rect 218 182 225 190
rect 251 161 258 258
rect 315 220 322 258
rect 355 220 362 328
rect 396 220 403 328
rect 437 255 444 328
rect 437 248 451 255
rect 437 225 451 232
rect 437 220 444 225
rect 495 220 502 516
rect 527 486 534 539
rect 527 366 534 438
rect 527 288 534 328
rect 251 110 258 131
rect 315 127 322 190
rect 355 128 362 190
rect 396 161 403 190
rect 437 161 444 190
rect 495 180 502 190
rect 495 142 502 150
rect 527 142 534 258
rect 563 227 570 564
rect 553 220 570 227
rect 560 190 567 195
rect 553 188 567 190
rect 560 180 567 188
rect 560 142 567 150
rect 396 120 403 131
rect 437 120 444 131
<< ndiffusion >>
rect 27 317 29 347
rect 36 317 38 347
rect 54 317 59 347
rect 66 317 88 347
rect 95 317 97 347
rect 113 317 115 347
rect 122 317 124 347
rect 27 252 29 282
rect 36 252 38 282
rect 144 252 146 282
rect 153 252 155 282
rect 310 328 315 366
rect 322 328 355 366
rect 362 328 369 366
rect 385 328 396 366
rect 403 328 437 366
rect 444 328 449 366
rect 246 258 251 288
rect 258 258 315 288
rect 322 258 333 288
rect 216 190 218 220
rect 225 190 230 220
rect 525 258 527 288
rect 534 258 540 288
rect 313 190 315 220
rect 322 190 355 220
rect 362 190 365 220
rect 429 190 437 220
rect 444 190 495 220
rect 502 190 506 220
rect 246 131 251 161
rect 258 131 263 161
rect 394 131 396 161
rect 403 131 437 161
rect 444 131 448 161
rect 557 150 560 180
rect 567 150 570 180
<< pdiffusion >>
rect 27 643 29 691
rect 36 643 38 691
rect 54 643 59 691
rect 66 643 68 691
rect 84 643 88 691
rect 95 643 97 691
rect 113 643 115 691
rect 122 643 125 691
rect 141 643 146 691
rect 153 643 156 691
rect 249 643 251 691
rect 258 643 260 691
rect 276 643 281 691
rect 288 643 290 691
rect 27 564 29 612
rect 36 564 38 612
rect 215 562 218 610
rect 225 562 230 610
rect 420 643 437 691
rect 444 643 454 691
rect 470 643 495 691
rect 502 643 505 691
rect 279 564 281 612
rect 288 564 316 612
rect 332 564 334 612
rect 341 564 351 612
rect 367 564 375 612
rect 382 564 384 612
rect 400 564 437 612
rect 444 564 446 612
rect 560 564 563 612
rect 570 564 580 612
rect 249 438 251 486
rect 258 438 261 486
rect 277 438 281 486
rect 288 438 290 486
rect 310 438 334 486
rect 341 438 349 486
rect 367 438 375 486
rect 382 438 384 486
rect 400 438 437 486
rect 444 438 447 486
rect 524 438 527 486
rect 534 438 540 486
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 188 86
rect 0 76 188 79
<< nohmic >>
rect 0 743 188 746
rect 0 736 8 743
rect 24 736 36 743
rect 52 736 64 743
rect 80 736 92 743
rect 108 736 120 743
rect 136 736 148 743
rect 164 736 188 743
<< ntransistor >>
rect 29 317 36 347
rect 59 317 66 347
rect 88 317 95 347
rect 115 317 122 347
rect 29 252 36 282
rect 146 252 153 282
rect 315 328 322 366
rect 355 328 362 366
rect 396 328 403 366
rect 437 328 444 366
rect 251 258 258 288
rect 315 258 322 288
rect 218 190 225 220
rect 527 258 534 288
rect 315 190 322 220
rect 355 190 362 220
rect 437 190 444 220
rect 495 190 502 220
rect 251 131 258 161
rect 396 131 403 161
rect 437 131 444 161
rect 560 150 567 180
<< ptransistor >>
rect 29 643 36 691
rect 59 643 66 691
rect 88 643 95 691
rect 115 643 122 691
rect 146 643 153 691
rect 251 643 258 691
rect 281 643 288 691
rect 29 564 36 612
rect 218 562 225 610
rect 437 643 444 691
rect 495 643 502 691
rect 281 564 288 612
rect 334 564 341 612
rect 375 564 382 612
rect 437 564 444 612
rect 563 564 570 612
rect 251 438 258 486
rect 281 438 288 486
rect 334 438 341 486
rect 375 438 382 486
rect 437 438 444 486
rect 527 438 534 486
<< polycontact >>
rect 316 695 332 711
rect 366 645 382 661
rect 59 583 75 599
rect 133 617 149 633
rect 116 575 132 591
rect 84 557 100 573
rect 132 377 148 393
rect 554 675 570 691
rect 518 539 534 555
rect 490 516 506 532
rect 209 372 225 388
rect 59 262 75 278
rect 37 226 53 242
rect 334 412 350 428
rect 437 412 453 428
rect 247 315 263 331
rect 439 232 455 248
rect 518 328 534 366
rect 387 190 403 220
rect 495 150 511 180
rect 544 190 560 220
rect 310 111 326 127
rect 351 111 368 128
<< ndiffcontact >>
rect 11 317 27 347
rect 38 317 54 347
rect 97 317 113 347
rect 124 317 140 347
rect 11 252 27 282
rect 38 252 54 282
rect 128 252 144 282
rect 155 252 171 282
rect 294 328 310 366
rect 369 328 385 366
rect 449 328 465 366
rect 230 258 246 288
rect 333 258 349 288
rect 200 190 216 220
rect 230 190 246 220
rect 509 258 525 288
rect 540 258 556 288
rect 297 190 313 220
rect 365 190 381 220
rect 413 190 429 220
rect 506 190 522 220
rect 230 131 246 161
rect 263 131 279 161
rect 378 131 394 161
rect 448 131 464 161
rect 541 150 557 180
rect 570 150 586 180
<< pdiffcontact >>
rect 11 643 27 691
rect 38 643 54 691
rect 68 643 84 691
rect 97 643 113 691
rect 125 643 141 691
rect 156 643 172 691
rect 233 643 249 691
rect 260 643 276 691
rect 290 643 306 691
rect 11 564 27 612
rect 38 564 54 612
rect 199 562 215 610
rect 230 562 246 610
rect 404 643 420 691
rect 454 643 470 691
rect 505 643 521 691
rect 263 564 279 612
rect 316 564 332 612
rect 351 564 367 612
rect 384 564 400 612
rect 446 564 462 612
rect 544 564 560 612
rect 580 564 596 612
rect 233 438 249 486
rect 261 438 277 486
rect 290 438 310 486
rect 349 438 367 486
rect 384 438 400 486
rect 447 438 463 486
rect 508 438 524 486
rect 540 438 557 486
<< psubstratetap >>
rect 6 79 22 95
rect 34 79 50 95
rect 62 79 78 95
rect 90 79 106 95
rect 118 79 134 95
rect 146 79 162 95
rect 404 80 421 97
<< nsubstratetap >>
rect 8 727 24 743
rect 36 727 52 743
rect 64 727 80 743
rect 92 727 108 743
rect 120 727 136 743
rect 148 727 164 743
rect 414 727 431 744
<< metal1 >>
rect 0 782 603 792
rect 0 759 118 769
rect 188 759 493 769
rect 509 759 603 769
rect 0 744 603 746
rect 0 743 414 744
rect 0 727 8 743
rect 24 727 36 743
rect 52 727 64 743
rect 80 727 92 743
rect 108 727 120 743
rect 136 727 148 743
rect 164 727 414 743
rect 431 727 603 744
rect 0 721 603 727
rect 11 691 27 721
rect 41 701 110 711
rect 41 691 51 701
rect 100 691 110 701
rect 125 691 141 721
rect 11 612 27 643
rect 71 629 81 643
rect 71 619 133 629
rect 54 583 59 599
rect 41 380 132 390
rect 41 347 51 380
rect 159 385 169 643
rect 199 634 215 721
rect 233 691 249 721
rect 260 701 316 711
rect 260 691 276 701
rect 454 701 554 711
rect 454 691 470 701
rect 554 691 570 695
rect 199 633 216 634
rect 290 633 306 643
rect 199 621 306 633
rect 316 645 366 655
rect 199 610 215 621
rect 263 612 279 621
rect 199 511 215 562
rect 316 612 332 645
rect 404 633 420 643
rect 505 633 521 643
rect 580 633 596 721
rect 351 623 596 633
rect 351 612 367 623
rect 446 612 462 623
rect 580 612 596 623
rect 230 549 246 562
rect 316 549 332 564
rect 230 539 332 549
rect 384 554 400 564
rect 384 544 518 554
rect 290 516 464 526
rect 480 516 490 526
rect 544 526 560 564
rect 506 516 560 526
rect 199 501 277 511
rect 261 486 277 501
rect 290 486 310 516
rect 580 506 596 564
rect 349 496 463 506
rect 349 486 367 496
rect 447 486 463 496
rect 508 496 596 506
rect 508 486 524 496
rect 463 438 508 486
rect 233 428 249 438
rect 384 428 400 438
rect 540 428 557 438
rect 233 418 334 428
rect 350 418 400 428
rect 453 418 557 428
rect 248 390 385 402
rect 159 375 209 385
rect 73 357 137 367
rect 14 307 24 317
rect 73 307 83 357
rect 127 347 137 357
rect 14 297 83 307
rect 54 262 59 278
rect 11 101 27 252
rect 97 101 113 317
rect 159 282 169 375
rect 248 353 261 390
rect 369 366 385 390
rect 200 341 261 353
rect 200 288 216 341
rect 247 314 263 315
rect 465 328 518 366
rect 294 318 310 328
rect 294 308 586 318
rect 200 258 230 288
rect 349 278 509 288
rect 128 101 144 252
rect 200 220 216 258
rect 230 247 246 258
rect 540 248 556 258
rect 230 235 429 247
rect 413 220 429 235
rect 455 232 556 248
rect 246 190 297 220
rect 381 190 387 220
rect 522 190 544 220
rect 200 161 216 190
rect 570 180 586 308
rect 200 131 230 161
rect 279 151 378 161
rect 511 150 541 180
rect 200 101 218 131
rect 309 111 310 127
rect 448 121 464 131
rect 368 111 464 121
rect 0 97 603 101
rect 0 95 404 97
rect 0 79 6 95
rect 22 79 34 95
rect 50 79 62 95
rect 78 79 90 95
rect 106 79 118 95
rect 134 79 146 95
rect 162 80 404 95
rect 421 80 603 97
rect 162 79 603 80
rect 0 76 603 79
rect 0 53 247 63
rect 263 53 603 63
rect 0 30 39 40
rect 53 30 603 40
rect 0 7 293 17
rect 309 7 603 17
<< m2contact >>
rect 118 757 132 771
rect 493 756 509 772
rect 118 591 132 605
rect 85 543 99 557
rect 554 695 570 711
rect 464 516 480 532
rect 39 212 53 226
rect 247 298 263 314
rect 293 111 309 127
rect 247 50 263 66
rect 39 28 53 42
rect 293 3 309 19
<< metal2 >>
rect 96 557 108 799
rect 119 605 131 757
rect 99 543 108 557
rect 40 42 52 212
rect 96 0 108 543
rect 466 532 478 799
rect 495 772 507 799
rect 495 711 507 756
rect 495 695 554 711
rect 247 66 263 298
rect 293 19 309 111
rect 466 0 478 516
rect 495 0 507 695
<< labels >>
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal2 96 799 108 799 5 D
rlabel metal1 0 76 0 101 1 GND!
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 3 Clock
rlabel metal2 96 0 108 0 1 D
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 603 7 603 17 7 nReset
rlabel metal1 603 30 603 40 7 Test
rlabel metal1 603 53 603 63 7 Clock
rlabel metal1 603 76 603 101 7 GND!
rlabel metal2 495 0 507 0 1 Q
rlabel metal2 466 0 478 0 1 nQ
rlabel metal1 603 759 603 769 7 Q
rlabel metal1 603 782 603 792 7 ScanReturn
rlabel metal2 495 799 507 799 5 Q
rlabel metal2 466 799 478 799 5 nQ
<< end >>
