magic
tech c035u
timestamp 1386362200
<< error_ps >>
rect 407 834 408 835
<< metal1 >>
rect 325 860 431 870
rect 205 836 407 846
rect 85 813 384 823
rect 469 813 504 823
rect 518 813 623 823
<< m2contact >>
rect 311 860 325 874
rect 431 858 445 872
rect 191 834 205 848
rect 407 834 421 848
rect 71 809 85 823
rect 384 811 398 825
rect 455 809 469 823
rect 504 811 518 825
rect 623 811 637 825
<< metal2 >>
rect 24 799 36 891
rect 72 799 84 809
rect 144 799 156 891
rect 192 799 204 834
rect 264 799 276 891
rect 312 799 324 860
rect 384 825 396 891
rect 408 848 420 891
rect 432 872 444 891
rect 384 799 396 811
rect 408 799 420 834
rect 432 799 444 858
rect 456 823 468 891
rect 456 799 468 809
rect 504 799 516 811
rect 552 799 564 891
rect 624 799 636 811
rect 672 799 684 891
use inv inv_2
timestamp 1386238110
transform 1 0 0 0 1 0
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 120 0 1 0
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 240 0 1 0
box 0 0 120 799
use nand3 nand3_0
timestamp 1386234893
transform 1 0 360 0 1 0
box 0 0 120 799
use inv inv_0
timestamp 1386238110
transform 1 0 480 0 1 0
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 600 0 1 0
box 0 0 120 799
<< labels >>
rlabel metal2 672 891 684 891 5 n2
rlabel metal2 552 891 564 891 5 n1
rlabel metal2 456 891 468 891 5 Y
rlabel metal2 432 891 444 891 5 C
rlabel metal2 408 891 420 891 5 B
rlabel metal2 384 891 396 891 5 A
rlabel metal2 24 891 36 891 5 NA
rlabel metal2 144 891 156 891 5 NB
rlabel metal2 264 891 276 891 5 NC
<< end >>
