magic
tech c035u
timestamp 1385631458
<< nwell >>
rect 2 597 122 746
rect 0 534 122 597
<< polysilicon >>
rect 30 597 37 605
rect 57 597 64 605
rect 84 597 91 605
rect 30 389 37 549
rect 57 451 64 549
rect 63 435 64 451
rect 30 363 37 373
rect 57 363 64 435
rect 84 416 91 549
rect 90 400 91 416
rect 83 386 91 400
rect 84 363 91 386
rect 30 325 37 333
rect 57 325 64 333
rect 84 325 91 333
<< ndiffusion >>
rect 28 333 30 363
rect 37 333 57 363
rect 64 333 84 363
rect 91 333 93 363
<< pdiffusion >>
rect 28 549 30 597
rect 37 549 39 597
rect 55 549 57 597
rect 64 549 66 597
rect 82 549 84 597
rect 91 549 93 597
<< pohmic >>
rect 2 79 8 86
rect 24 79 36 86
rect 52 79 92 86
rect 108 79 122 86
rect 2 76 122 79
<< nohmic >>
rect 2 743 119 746
rect 2 736 8 743
rect 24 736 36 743
rect 52 736 64 743
rect 80 736 119 743
<< ntransistor >>
rect 30 333 37 363
rect 57 333 64 363
rect 84 333 91 363
<< ptransistor >>
rect 30 549 37 597
rect 57 549 64 597
rect 84 549 91 597
<< polycontact >>
rect 47 435 63 451
rect 26 373 42 389
rect 74 400 90 416
<< ndiffcontact >>
rect 12 333 28 363
rect 93 333 109 363
<< pdiffcontact >>
rect 12 549 28 597
rect 39 549 55 597
rect 66 549 82 597
rect 93 549 109 597
<< psubstratetap >>
rect 8 79 24 95
rect 36 79 52 95
rect 92 79 108 95
<< nsubstratetap >>
rect 8 727 24 743
rect 36 727 52 743
rect 64 727 80 743
<< metal1 >>
rect 2 782 122 792
rect 2 759 122 769
rect 2 743 122 746
rect 2 727 8 743
rect 24 727 36 743
rect 52 727 64 743
rect 80 727 122 743
rect 2 721 122 727
rect 12 597 28 721
rect 66 597 82 721
rect 45 499 55 549
rect 99 499 109 549
rect 45 489 99 499
rect 100 363 110 485
rect 109 333 110 363
rect 12 101 28 333
rect 2 95 122 101
rect 2 79 8 95
rect 24 79 36 95
rect 52 79 92 95
rect 108 79 122 95
rect 2 76 122 79
rect 2 53 122 63
rect 2 30 122 40
rect 2 7 122 17
<< m2contact >>
rect 99 485 113 499
rect 48 421 62 435
rect 26 389 40 403
rect 74 386 88 400
<< metal2 >>
rect 26 597 38 799
rect 26 549 39 597
rect 26 403 38 549
rect 50 451 62 799
rect 50 435 63 451
rect 26 373 40 389
rect 26 0 38 373
rect 50 0 62 421
rect 74 416 86 799
rect 98 499 110 799
rect 98 485 99 499
rect 74 400 87 416
rect 74 0 86 386
rect 98 0 110 485
<< labels >>
rlabel metal1 2 77 2 101 3 GND!
rlabel metal1 2 7 2 17 2 nReset
rlabel metal1 2 30 2 40 3 Test
rlabel metal1 2 53 2 63 3 Clock
rlabel metal1 122 77 122 101 7 GND!
rlabel metal1 122 7 122 17 8 nReset
rlabel metal1 122 30 122 40 7 Test
rlabel metal1 122 53 122 63 7 Clock
rlabel metal2 98 0 110 0 1 Y
rlabel metal2 74 0 86 0 1 C
rlabel metal2 26 0 38 0 1 A
rlabel metal2 50 0 62 0 1 B
rlabel metal2 98 799 110 799 5 Y
rlabel metal2 74 799 86 799 5 C
rlabel metal2 50 799 62 799 5 B
rlabel metal2 26 799 38 799 5 A
rlabel metal1 122 782 122 792 6 ScanReturn
rlabel metal1 122 759 122 769 7 Scan
rlabel metal1 122 721 122 746 7 Vdd!
rlabel metal1 2 782 2 792 4 ScanReturn
rlabel metal1 2 759 2 769 3 Scan
rlabel metal1 2 721 2 746 3 Vdd!
<< end >>
