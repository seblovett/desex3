magic
tech c035u
timestamp 1385125399
<< metal1 >>
rect 0 745 10 770
rect 0 110 10 135
<< metal2 >>
rect 34 0 46 37
rect 58 0 70 37
rect 82 27 94 37
rect 154 27 166 37
rect 274 27 286 37
rect 82 15 286 27
rect 82 0 94 15
use nor2 nor2_0
timestamp 1385124540
transform 1 0 10 0 1 37
box 0 0 120 783
use inv inv_0
timestamp 1385124685
transform 1 0 130 0 1 37
box 0 0 120 783
use inv inv_1
timestamp 1385124685
transform 1 0 250 0 1 37
box 0 0 120 783
<< labels >>
rlabel metal2 34 0 46 0 1 A
rlabel metal2 58 0 70 0 1 B
rlabel metal2 82 0 94 0 1 Y
rlabel metal1 0 110 0 135 3 GND!
rlabel metal1 0 745 0 770 3 Vdd!
<< end >>
