magic
tech c035u
timestamp 1385034376
<< nwell >>
rect 202 524 1499 736
rect 202 489 1387 524
rect 202 488 1371 489
rect 324 396 641 488
rect 689 396 1006 488
rect 1054 396 1371 488
rect 377 395 423 396
rect 742 395 788 396
rect 1107 395 1153 396
<< polysilicon >>
rect 535 686 542 694
rect 562 686 569 694
rect 589 686 596 694
rect 616 686 623 694
rect 900 686 907 694
rect 927 686 934 694
rect 954 686 961 694
rect 981 686 988 694
rect 1265 686 1272 694
rect 1292 686 1299 694
rect 1319 686 1326 694
rect 1346 686 1353 694
rect 452 608 459 616
rect 479 608 486 616
rect 397 553 404 561
rect 342 454 349 462
rect 817 608 824 616
rect 844 608 851 616
rect 762 553 769 561
rect 707 454 714 462
rect 1182 608 1189 616
rect 1209 608 1216 616
rect 1127 553 1134 561
rect 1072 454 1079 462
rect 1451 637 1453 653
rect 1446 592 1453 637
rect 1446 496 1453 544
rect 1446 458 1453 466
rect 342 382 349 396
rect 397 382 404 396
rect 452 383 459 396
rect 347 366 349 382
rect 402 366 404 382
rect 457 379 459 383
rect 479 379 486 396
rect 535 383 542 396
rect 457 372 486 379
rect 457 367 459 372
rect 540 379 542 383
rect 562 379 569 396
rect 589 379 596 396
rect 616 379 623 396
rect 707 382 714 396
rect 762 382 769 396
rect 817 383 824 396
rect 540 372 623 379
rect 540 367 542 372
rect 342 356 349 366
rect 397 356 404 366
rect 452 356 459 367
rect 535 356 542 367
rect 562 356 569 372
rect 712 366 714 382
rect 767 366 769 382
rect 822 379 824 383
rect 844 379 851 396
rect 900 383 907 396
rect 822 372 851 379
rect 822 367 824 372
rect 905 379 907 383
rect 927 379 934 396
rect 954 379 961 396
rect 981 379 988 396
rect 1072 382 1079 396
rect 1127 382 1134 396
rect 1182 383 1189 396
rect 905 372 988 379
rect 905 367 907 372
rect 707 356 714 366
rect 762 356 769 366
rect 817 356 824 367
rect 900 356 907 367
rect 927 356 934 372
rect 1077 366 1079 382
rect 1132 366 1134 382
rect 1187 379 1189 383
rect 1209 379 1216 396
rect 1265 383 1272 396
rect 1187 372 1216 379
rect 1187 367 1189 372
rect 1270 379 1272 383
rect 1292 379 1299 396
rect 1319 379 1326 396
rect 1346 379 1353 396
rect 1270 372 1353 379
rect 1270 367 1272 372
rect 1072 356 1079 366
rect 1127 356 1134 366
rect 1182 356 1189 367
rect 1265 356 1272 367
rect 1292 356 1299 372
rect 342 328 349 336
rect 397 294 404 302
rect 452 202 459 210
rect 707 328 714 336
rect 762 294 769 302
rect 817 202 824 210
rect 1072 328 1079 336
rect 1127 294 1134 302
rect 1182 202 1189 210
rect 535 148 542 156
rect 562 148 569 156
rect 900 148 907 156
rect 927 148 934 156
rect 1265 148 1272 156
rect 1292 148 1299 156
<< ndiffusion >>
rect 1444 466 1446 496
rect 1453 466 1455 496
rect 340 336 342 356
rect 349 336 351 356
rect 395 302 397 356
rect 404 302 406 356
rect 450 210 452 356
rect 459 210 461 356
rect 533 156 535 356
rect 542 156 544 356
rect 560 156 562 356
rect 569 156 571 356
rect 705 336 707 356
rect 714 336 716 356
rect 760 302 762 356
rect 769 302 771 356
rect 815 210 817 356
rect 824 210 826 356
rect 898 156 900 356
rect 907 156 909 356
rect 925 156 927 356
rect 934 156 936 356
rect 1070 336 1072 356
rect 1079 336 1081 356
rect 1125 302 1127 356
rect 1134 302 1136 356
rect 1180 210 1182 356
rect 1189 210 1191 356
rect 1263 156 1265 356
rect 1272 156 1274 356
rect 1290 156 1292 356
rect 1299 156 1301 356
<< pdiffusion >>
rect 340 396 342 454
rect 349 396 351 454
rect 395 396 397 553
rect 404 396 406 553
rect 450 396 452 608
rect 459 396 461 608
rect 477 396 479 608
rect 486 396 488 608
rect 533 396 535 686
rect 542 396 544 686
rect 560 396 562 686
rect 569 396 571 686
rect 587 396 589 686
rect 596 396 598 686
rect 614 396 616 686
rect 623 396 625 686
rect 705 396 707 454
rect 714 396 716 454
rect 760 396 762 553
rect 769 396 771 553
rect 815 396 817 608
rect 824 396 826 608
rect 842 396 844 608
rect 851 396 853 608
rect 898 396 900 686
rect 907 396 909 686
rect 925 396 927 686
rect 934 396 936 686
rect 952 396 954 686
rect 961 396 963 686
rect 979 396 981 686
rect 988 396 990 686
rect 1070 396 1072 454
rect 1079 396 1081 454
rect 1125 396 1127 553
rect 1134 396 1136 553
rect 1180 396 1182 608
rect 1189 396 1191 608
rect 1207 396 1209 608
rect 1216 396 1218 608
rect 1263 396 1265 686
rect 1272 396 1274 686
rect 1290 396 1292 686
rect 1299 396 1301 686
rect 1317 396 1319 686
rect 1326 396 1328 686
rect 1344 396 1346 686
rect 1353 396 1355 686
rect 1444 544 1446 592
rect 1453 544 1455 592
<< pohmic >>
rect 324 76 326 86
rect 342 76 354 86
rect 370 76 382 86
rect 398 76 410 86
rect 426 76 438 86
rect 454 76 466 86
rect 482 76 494 86
rect 510 76 522 86
rect 539 76 551 86
rect 567 76 579 86
rect 595 76 607 86
rect 623 76 635 86
rect 651 76 663 86
rect 679 76 691 86
rect 707 76 719 86
rect 735 76 747 86
rect 763 76 775 86
rect 791 76 803 86
rect 819 76 831 86
rect 847 76 859 86
rect 875 76 887 86
rect 904 76 916 86
rect 932 76 944 86
rect 960 76 972 86
rect 988 76 1000 86
rect 1016 76 1028 86
rect 1044 76 1056 86
rect 1072 76 1084 86
rect 1100 76 1112 86
rect 1128 76 1140 86
rect 1156 76 1168 86
rect 1184 76 1196 86
rect 1212 76 1224 86
rect 1240 76 1252 86
rect 1269 76 1281 86
rect 1297 76 1309 86
rect 1325 76 1337 86
rect 1353 76 1365 86
rect 1381 76 1393 86
rect 1409 76 1421 86
rect 1437 76 1449 86
rect 1465 76 1477 86
rect 1493 76 1499 86
<< nohmic >>
rect 202 726 214 736
rect 230 726 242 736
rect 258 726 270 736
rect 286 726 298 736
rect 314 726 326 736
rect 342 726 354 736
rect 370 726 382 736
rect 398 726 410 736
rect 426 726 438 736
rect 454 726 466 736
rect 482 726 494 736
rect 510 726 522 736
rect 539 726 551 736
rect 567 726 579 736
rect 595 726 607 736
rect 623 726 635 736
rect 651 726 663 736
rect 679 726 691 736
rect 707 726 719 736
rect 735 726 747 736
rect 763 726 775 736
rect 791 726 803 736
rect 819 726 831 736
rect 847 726 859 736
rect 875 726 887 736
rect 904 726 916 736
rect 932 726 944 736
rect 960 726 972 736
rect 988 726 1000 736
rect 1016 726 1028 736
rect 1044 726 1056 736
rect 1072 726 1084 736
rect 1100 726 1112 736
rect 1128 726 1140 736
rect 1156 726 1168 736
rect 1184 726 1196 736
rect 1212 726 1224 736
rect 1240 726 1252 736
rect 1269 726 1281 736
rect 1297 726 1309 736
rect 1325 726 1337 736
rect 1353 726 1365 736
rect 1381 726 1393 736
rect 1409 726 1421 736
rect 1437 726 1449 736
rect 1465 726 1477 736
rect 1493 726 1499 736
<< ntransistor >>
rect 1446 466 1453 496
rect 342 336 349 356
rect 397 302 404 356
rect 452 210 459 356
rect 535 156 542 356
rect 562 156 569 356
rect 707 336 714 356
rect 762 302 769 356
rect 817 210 824 356
rect 900 156 907 356
rect 927 156 934 356
rect 1072 336 1079 356
rect 1127 302 1134 356
rect 1182 210 1189 356
rect 1265 156 1272 356
rect 1292 156 1299 356
<< ptransistor >>
rect 342 396 349 454
rect 397 396 404 553
rect 452 396 459 608
rect 479 396 486 608
rect 535 396 542 686
rect 562 396 569 686
rect 589 396 596 686
rect 616 396 623 686
rect 707 396 714 454
rect 762 396 769 553
rect 817 396 824 608
rect 844 396 851 608
rect 900 396 907 686
rect 927 396 934 686
rect 954 396 961 686
rect 981 396 988 686
rect 1072 396 1079 454
rect 1127 396 1134 553
rect 1182 396 1189 608
rect 1209 396 1216 608
rect 1265 396 1272 686
rect 1292 396 1299 686
rect 1319 396 1326 686
rect 1346 396 1353 686
rect 1446 544 1453 592
<< polycontact >>
rect 1435 637 1451 653
rect 331 366 347 382
rect 386 366 402 382
rect 441 367 457 383
rect 524 367 540 383
rect 696 366 712 382
rect 751 366 767 382
rect 806 367 822 383
rect 889 367 905 383
rect 1061 366 1077 382
rect 1116 366 1132 382
rect 1171 367 1187 383
rect 1254 367 1270 383
<< ndiffcontact >>
rect 1428 466 1444 496
rect 1455 466 1471 496
rect 324 336 340 356
rect 351 336 367 356
rect 379 302 395 356
rect 406 302 422 356
rect 434 210 450 356
rect 461 210 477 356
rect 517 156 533 356
rect 544 156 560 356
rect 571 156 587 356
rect 689 336 705 356
rect 716 336 732 356
rect 744 302 760 356
rect 771 302 787 356
rect 799 210 815 356
rect 826 210 842 356
rect 882 156 898 356
rect 909 156 925 356
rect 936 156 952 356
rect 1054 336 1070 356
rect 1081 336 1097 356
rect 1109 302 1125 356
rect 1136 302 1152 356
rect 1164 210 1180 356
rect 1191 210 1207 356
rect 1247 156 1263 356
rect 1274 156 1290 356
rect 1301 156 1317 356
<< pdiffcontact >>
rect 324 396 340 454
rect 351 396 367 454
rect 379 396 395 553
rect 406 396 422 553
rect 434 396 450 608
rect 461 396 477 608
rect 488 396 504 608
rect 517 396 533 686
rect 544 396 560 686
rect 571 396 587 686
rect 598 396 614 686
rect 625 396 641 686
rect 689 396 705 454
rect 716 396 732 454
rect 744 396 760 553
rect 771 396 787 553
rect 799 396 815 608
rect 826 396 842 608
rect 853 396 869 608
rect 882 396 898 686
rect 909 396 925 686
rect 936 396 952 686
rect 963 396 979 686
rect 990 396 1006 686
rect 1054 396 1070 454
rect 1081 396 1097 454
rect 1109 396 1125 553
rect 1136 396 1152 553
rect 1164 396 1180 608
rect 1191 396 1207 608
rect 1218 396 1234 608
rect 1247 396 1263 686
rect 1274 396 1290 686
rect 1301 396 1317 686
rect 1328 396 1344 686
rect 1355 396 1371 686
rect 1428 544 1444 592
rect 1455 544 1471 592
<< psubstratetap >>
rect 326 76 342 92
rect 354 76 370 92
rect 382 76 398 92
rect 410 76 426 92
rect 438 76 454 92
rect 466 76 482 92
rect 494 76 510 92
rect 522 76 539 92
rect 551 76 567 92
rect 579 76 595 92
rect 607 76 623 92
rect 635 76 651 92
rect 663 76 679 92
rect 691 76 707 92
rect 719 76 735 92
rect 747 76 763 92
rect 775 76 791 92
rect 803 76 819 92
rect 831 76 847 92
rect 859 76 875 92
rect 887 76 904 92
rect 916 76 932 92
rect 944 76 960 92
rect 972 76 988 92
rect 1000 76 1016 92
rect 1028 76 1044 92
rect 1056 76 1072 92
rect 1084 76 1100 92
rect 1112 76 1128 92
rect 1140 76 1156 92
rect 1168 76 1184 92
rect 1196 76 1212 92
rect 1224 76 1240 92
rect 1252 76 1269 92
rect 1281 76 1297 92
rect 1309 76 1325 92
rect 1337 76 1353 92
rect 1365 76 1381 92
rect 1393 76 1409 92
rect 1421 76 1437 92
rect 1449 76 1465 92
rect 1477 76 1493 92
<< nsubstratetap >>
rect 214 720 230 736
rect 242 720 258 736
rect 270 720 286 736
rect 298 720 314 736
rect 326 720 342 736
rect 354 720 370 736
rect 382 720 398 736
rect 410 720 426 736
rect 438 720 454 736
rect 466 720 482 736
rect 494 720 510 736
rect 522 720 539 736
rect 551 720 567 736
rect 579 720 595 736
rect 607 720 623 736
rect 635 720 651 736
rect 663 720 679 736
rect 691 720 707 736
rect 719 720 735 736
rect 747 720 763 736
rect 775 720 791 736
rect 803 720 819 736
rect 831 720 847 736
rect 859 720 875 736
rect 887 720 904 736
rect 916 720 932 736
rect 944 720 960 736
rect 972 720 988 736
rect 1000 720 1016 736
rect 1028 720 1044 736
rect 1056 720 1072 736
rect 1084 720 1100 736
rect 1112 720 1128 736
rect 1140 720 1156 736
rect 1168 720 1184 736
rect 1196 720 1212 736
rect 1224 720 1240 736
rect 1252 720 1269 736
rect 1281 720 1297 736
rect 1309 720 1325 736
rect 1337 720 1353 736
rect 1365 720 1381 736
rect 1393 720 1409 736
rect 1421 720 1437 736
rect 1449 720 1465 736
rect 1477 720 1493 736
<< metal1 >>
rect 236 772 1413 782
rect 1457 772 1499 782
rect 236 749 1499 759
rect 200 720 214 736
rect 230 720 242 736
rect 258 720 270 736
rect 286 720 298 736
rect 314 720 326 736
rect 342 720 354 736
rect 370 720 382 736
rect 398 720 410 736
rect 426 720 438 736
rect 454 720 466 736
rect 482 720 494 736
rect 510 720 522 736
rect 539 720 551 736
rect 567 720 579 736
rect 595 720 607 736
rect 623 720 635 736
rect 651 720 663 736
rect 679 720 691 736
rect 707 720 719 736
rect 735 720 747 736
rect 763 720 775 736
rect 791 720 803 736
rect 819 720 831 736
rect 847 720 859 736
rect 875 720 887 736
rect 904 720 916 736
rect 932 720 944 736
rect 960 720 972 736
rect 988 720 1000 736
rect 1016 720 1028 736
rect 1044 720 1056 736
rect 1072 720 1084 736
rect 1100 720 1112 736
rect 1128 720 1140 736
rect 1156 720 1168 736
rect 1184 720 1196 736
rect 1212 720 1224 736
rect 1240 720 1252 736
rect 1269 720 1281 736
rect 1297 720 1309 736
rect 1325 720 1337 736
rect 1353 720 1365 736
rect 1381 720 1393 736
rect 1409 720 1421 736
rect 1437 720 1449 736
rect 1465 720 1477 736
rect 1493 720 1499 736
rect 200 711 1499 720
rect 324 454 340 711
rect 379 553 395 711
rect 434 608 450 711
rect 488 608 504 711
rect 517 686 533 711
rect 571 686 587 711
rect 625 686 641 711
rect 689 454 705 711
rect 744 553 760 711
rect 799 608 815 711
rect 853 608 869 711
rect 882 686 898 711
rect 936 686 952 711
rect 990 686 1006 711
rect 1054 454 1070 711
rect 1109 553 1125 711
rect 1164 608 1180 711
rect 1218 608 1234 711
rect 1247 686 1263 711
rect 1301 686 1317 711
rect 1355 686 1371 711
rect 1437 653 1451 659
rect 1461 592 1471 711
rect 1428 496 1438 544
rect 284 369 331 379
rect 357 379 367 396
rect 357 369 386 379
rect 357 356 367 369
rect 412 380 422 396
rect 412 370 441 380
rect 412 356 422 370
rect 467 380 477 396
rect 467 370 524 380
rect 467 356 477 370
rect 550 381 560 396
rect 604 383 614 396
rect 550 371 602 381
rect 550 356 560 371
rect 685 369 696 379
rect 722 379 732 396
rect 722 369 751 379
rect 722 356 732 369
rect 777 380 787 396
rect 777 370 806 380
rect 777 356 787 370
rect 832 380 842 396
rect 832 370 889 380
rect 832 356 842 370
rect 915 381 925 396
rect 969 383 979 396
rect 915 371 965 381
rect 915 356 925 371
rect 1051 369 1061 379
rect 1087 379 1097 396
rect 1087 369 1116 379
rect 1087 356 1097 369
rect 1142 380 1152 396
rect 1142 370 1171 380
rect 1142 356 1152 370
rect 1197 380 1207 396
rect 1197 370 1254 380
rect 1197 356 1207 370
rect 1280 381 1290 396
rect 1334 383 1344 396
rect 1280 371 1328 381
rect 1280 356 1290 371
rect 1342 381 1344 383
rect 1342 371 1387 381
rect 324 101 340 336
rect 379 101 395 302
rect 434 101 450 210
rect 517 101 533 156
rect 571 101 587 156
rect 689 101 705 336
rect 744 101 760 302
rect 799 101 815 210
rect 882 101 898 156
rect 936 101 952 156
rect 1054 101 1070 336
rect 1109 101 1125 302
rect 1164 101 1180 210
rect 1247 101 1263 156
rect 1301 101 1317 156
rect 1455 101 1465 466
rect 324 92 1499 101
rect 324 76 326 92
rect 342 76 354 92
rect 370 76 382 92
rect 398 76 410 92
rect 426 76 438 92
rect 454 76 466 92
rect 482 76 494 92
rect 510 76 522 92
rect 539 76 551 92
rect 567 76 579 92
rect 595 76 607 92
rect 623 76 635 92
rect 651 76 663 92
rect 679 76 691 92
rect 707 76 719 92
rect 735 76 747 92
rect 763 76 775 92
rect 791 76 803 92
rect 819 76 831 92
rect 847 76 859 92
rect 875 76 887 92
rect 904 76 916 92
rect 932 76 944 92
rect 960 76 972 92
rect 988 76 1000 92
rect 1016 76 1028 92
rect 1044 76 1056 92
rect 1072 76 1084 92
rect 1100 76 1112 92
rect 1128 76 1140 92
rect 1156 76 1168 92
rect 1184 76 1196 92
rect 1212 76 1224 92
rect 1240 76 1252 92
rect 1269 76 1281 92
rect 1297 76 1309 92
rect 1325 76 1337 92
rect 1353 76 1365 92
rect 1381 76 1393 92
rect 1409 76 1421 92
rect 1437 76 1449 92
rect 1465 76 1477 92
rect 1493 76 1499 92
rect 617 53 1499 63
rect 260 30 671 40
rect 980 30 1499 40
rect 308 7 1036 17
rect 1343 7 1499 17
<< m2contact >>
rect 222 771 236 785
rect 1413 771 1427 785
rect 1443 771 1457 785
rect 222 747 236 761
rect 0 711 200 736
rect 1437 659 1451 673
rect 1414 578 1428 592
rect 270 367 284 381
rect 602 369 616 383
rect 671 367 685 381
rect 965 369 979 383
rect 1037 367 1051 381
rect 1328 369 1342 383
rect 603 51 617 65
rect 246 29 260 43
rect 671 28 685 42
rect 966 28 980 42
rect 294 5 308 19
rect 1036 5 1050 19
rect 1329 5 1343 19
<< metal2 >>
rect 0 736 200 790
rect 223 785 235 790
rect 0 0 200 711
rect 223 0 235 747
rect 247 43 259 790
rect 271 381 283 790
rect 247 0 259 29
rect 271 0 283 367
rect 295 19 307 790
rect 1415 592 1427 771
rect 1443 673 1455 771
rect 1451 659 1455 673
rect 604 65 616 369
rect 672 42 684 367
rect 967 42 979 369
rect 1037 19 1049 367
rect 1330 19 1342 369
rect 295 0 307 5
<< labels >>
rlabel metal1 1499 772 1499 782 7 nSDO
rlabel metal1 1499 749 1499 759 7 SDI
rlabel metal1 1499 711 1499 736 7 Vdd!
rlabel metal1 1499 76 1499 101 7 GND!
rlabel metal1 1499 53 1499 63 7 ClockOut
rlabel metal1 1499 30 1499 40 7 TestOut
rlabel metal1 1499 7 1499 17 7 nResetOut
rlabel metal2 247 0 259 0 1 Test
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 295 0 307 0 1 nReset
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 295 790 307 790 5 nReset
rlabel metal2 271 790 283 790 5 Clock
rlabel metal2 247 790 259 790 5 Test
rlabel metal2 223 790 235 790 5 SDO
rlabel metal2 0 790 200 790 5 Vdd!
<< end >>
