magic
tech c035u
timestamp 1385751497
<< nwell >>
rect 202 490 1464 736
rect 202 488 644 490
rect 352 398 644 488
rect 689 398 981 490
rect 1026 398 1464 490
rect 405 397 451 398
rect 742 397 788 398
rect 1079 397 1125 398
rect 1318 392 1464 398
<< polysilicon >>
rect 538 688 545 696
rect 565 688 572 696
rect 592 688 599 696
rect 619 688 626 696
rect 875 688 882 696
rect 902 688 909 696
rect 929 688 936 696
rect 956 688 963 696
rect 1212 688 1219 696
rect 1239 688 1246 696
rect 1266 688 1273 696
rect 1293 688 1300 696
rect 480 610 487 618
rect 507 610 514 618
rect 425 555 432 563
rect 370 456 377 464
rect 817 610 824 618
rect 844 610 851 618
rect 762 555 769 563
rect 707 456 714 464
rect 1154 610 1161 618
rect 1181 610 1188 618
rect 1099 555 1106 563
rect 1044 456 1051 464
rect 1394 506 1396 522
rect 1389 461 1396 506
rect 370 384 377 398
rect 425 384 432 398
rect 480 385 487 398
rect 375 368 377 384
rect 430 368 432 384
rect 485 381 487 385
rect 507 381 514 398
rect 538 385 545 398
rect 485 374 514 381
rect 485 369 487 374
rect 543 381 545 385
rect 565 381 572 398
rect 592 381 599 398
rect 619 381 626 398
rect 707 384 714 398
rect 762 384 769 398
rect 817 385 824 398
rect 543 374 626 381
rect 543 369 545 374
rect 370 358 377 368
rect 425 358 432 368
rect 480 358 487 369
rect 538 358 545 369
rect 565 358 572 374
rect 712 368 714 384
rect 767 368 769 384
rect 822 381 824 385
rect 844 381 851 398
rect 875 385 882 398
rect 822 374 851 381
rect 822 369 824 374
rect 880 381 882 385
rect 902 381 909 398
rect 929 381 936 398
rect 956 381 963 398
rect 1044 384 1051 398
rect 1099 384 1106 398
rect 1154 385 1161 398
rect 880 374 963 381
rect 880 369 882 374
rect 707 358 714 368
rect 762 358 769 368
rect 817 358 824 369
rect 875 358 882 369
rect 902 358 909 374
rect 1049 368 1051 384
rect 1104 368 1106 384
rect 1159 381 1161 385
rect 1181 381 1188 398
rect 1212 385 1219 398
rect 1159 374 1188 381
rect 1159 369 1161 374
rect 1217 381 1219 385
rect 1239 381 1246 398
rect 1266 381 1273 398
rect 1293 381 1300 398
rect 1217 374 1300 381
rect 1217 369 1219 374
rect 1044 358 1051 368
rect 1099 358 1106 368
rect 1154 358 1161 369
rect 1212 358 1219 369
rect 1239 358 1246 374
rect 1389 367 1396 413
rect 370 330 377 338
rect 425 296 432 304
rect 480 204 487 212
rect 707 330 714 338
rect 762 296 769 304
rect 817 204 824 212
rect 1044 330 1051 338
rect 1099 296 1106 304
rect 1154 204 1161 212
rect 1389 329 1396 337
rect 538 150 545 158
rect 565 150 572 158
rect 875 150 882 158
rect 902 150 909 158
rect 1212 150 1219 158
rect 1239 150 1246 158
<< ndiffusion >>
rect 368 338 370 358
rect 377 338 379 358
rect 423 304 425 358
rect 432 304 434 358
rect 478 212 480 358
rect 487 212 489 358
rect 536 158 538 358
rect 545 158 547 358
rect 563 158 565 358
rect 572 158 574 358
rect 705 338 707 358
rect 714 338 716 358
rect 760 304 762 358
rect 769 304 771 358
rect 815 212 817 358
rect 824 212 826 358
rect 873 158 875 358
rect 882 158 884 358
rect 900 158 902 358
rect 909 158 911 358
rect 1042 338 1044 358
rect 1051 338 1053 358
rect 1097 304 1099 358
rect 1106 304 1108 358
rect 1152 212 1154 358
rect 1161 212 1163 358
rect 1210 158 1212 358
rect 1219 158 1221 358
rect 1237 158 1239 358
rect 1246 158 1248 358
rect 1387 337 1389 367
rect 1396 337 1398 367
<< pdiffusion >>
rect 368 398 370 456
rect 377 398 379 456
rect 423 398 425 555
rect 432 398 434 555
rect 478 398 480 610
rect 487 398 489 610
rect 505 398 507 610
rect 514 398 516 610
rect 536 398 538 688
rect 545 398 547 688
rect 563 398 565 688
rect 572 398 574 688
rect 590 398 592 688
rect 599 398 601 688
rect 617 398 619 688
rect 626 398 628 688
rect 705 398 707 456
rect 714 398 716 456
rect 760 398 762 555
rect 769 398 771 555
rect 815 398 817 610
rect 824 398 826 610
rect 842 398 844 610
rect 851 398 853 610
rect 873 398 875 688
rect 882 398 884 688
rect 900 398 902 688
rect 909 398 911 688
rect 927 398 929 688
rect 936 398 938 688
rect 954 398 956 688
rect 963 398 965 688
rect 1042 398 1044 456
rect 1051 398 1053 456
rect 1097 398 1099 555
rect 1106 398 1108 555
rect 1152 398 1154 610
rect 1161 398 1163 610
rect 1179 398 1181 610
rect 1188 398 1190 610
rect 1210 398 1212 688
rect 1219 398 1221 688
rect 1237 398 1239 688
rect 1246 398 1248 688
rect 1264 398 1266 688
rect 1273 398 1275 688
rect 1291 398 1293 688
rect 1300 398 1302 688
rect 1387 413 1389 461
rect 1396 413 1398 461
<< pohmic >>
rect 320 66 326 76
rect 342 66 354 76
rect 370 66 382 76
rect 398 66 410 76
rect 426 66 438 76
rect 454 66 466 76
rect 482 66 494 76
rect 510 66 522 76
rect 538 66 550 76
rect 567 66 579 76
rect 595 66 607 76
rect 623 66 635 76
rect 651 66 663 76
rect 679 66 691 76
rect 707 66 719 76
rect 735 66 747 76
rect 763 66 775 76
rect 791 66 803 76
rect 819 66 831 76
rect 847 66 859 76
rect 875 66 887 76
rect 904 66 916 76
rect 932 66 944 76
rect 960 66 972 76
rect 988 66 1000 76
rect 1016 66 1028 76
rect 1044 66 1056 76
rect 1072 66 1084 76
rect 1100 66 1112 76
rect 1128 66 1140 76
rect 1156 66 1168 76
rect 1184 66 1196 76
rect 1212 66 1224 76
rect 1241 66 1253 76
rect 1269 66 1281 76
rect 1297 66 1309 76
rect 1325 66 1337 76
rect 1353 66 1365 76
rect 1381 66 1393 76
rect 1409 66 1421 76
rect 1437 66 1464 76
<< nohmic >>
rect 202 726 214 736
rect 230 726 242 736
rect 258 726 270 736
rect 286 726 298 736
rect 314 726 326 736
rect 342 726 354 736
rect 370 726 382 736
rect 398 726 410 736
rect 426 726 438 736
rect 454 726 466 736
rect 482 726 494 736
rect 510 726 522 736
rect 538 726 550 736
rect 567 726 579 736
rect 595 726 607 736
rect 623 726 635 736
rect 651 726 663 736
rect 679 726 691 736
rect 707 726 719 736
rect 735 726 747 736
rect 763 726 775 736
rect 791 726 803 736
rect 819 726 831 736
rect 847 726 859 736
rect 875 726 887 736
rect 904 726 916 736
rect 932 726 944 736
rect 960 726 972 736
rect 988 726 1000 736
rect 1016 726 1028 736
rect 1044 726 1056 736
rect 1072 726 1084 736
rect 1100 726 1112 736
rect 1128 726 1140 736
rect 1156 726 1168 736
rect 1184 726 1196 736
rect 1212 726 1224 736
rect 1241 726 1253 736
rect 1269 726 1281 736
rect 1297 726 1309 736
rect 1325 726 1337 736
rect 1353 726 1365 736
rect 1381 726 1393 736
rect 1409 726 1421 736
rect 1437 726 1464 736
<< ntransistor >>
rect 370 338 377 358
rect 425 304 432 358
rect 480 212 487 358
rect 538 158 545 358
rect 565 158 572 358
rect 707 338 714 358
rect 762 304 769 358
rect 817 212 824 358
rect 875 158 882 358
rect 902 158 909 358
rect 1044 338 1051 358
rect 1099 304 1106 358
rect 1154 212 1161 358
rect 1212 158 1219 358
rect 1239 158 1246 358
rect 1389 337 1396 367
<< ptransistor >>
rect 370 398 377 456
rect 425 398 432 555
rect 480 398 487 610
rect 507 398 514 610
rect 538 398 545 688
rect 565 398 572 688
rect 592 398 599 688
rect 619 398 626 688
rect 707 398 714 456
rect 762 398 769 555
rect 817 398 824 610
rect 844 398 851 610
rect 875 398 882 688
rect 902 398 909 688
rect 929 398 936 688
rect 956 398 963 688
rect 1044 398 1051 456
rect 1099 398 1106 555
rect 1154 398 1161 610
rect 1181 398 1188 610
rect 1212 398 1219 688
rect 1239 398 1246 688
rect 1266 398 1273 688
rect 1293 398 1300 688
rect 1389 413 1396 461
<< polycontact >>
rect 1378 506 1394 522
rect 359 368 375 384
rect 414 368 430 384
rect 469 369 485 385
rect 527 369 543 385
rect 696 368 712 384
rect 751 368 767 384
rect 806 369 822 385
rect 864 369 880 385
rect 1033 368 1049 384
rect 1088 368 1104 384
rect 1143 369 1159 385
rect 1201 369 1217 385
<< ndiffcontact >>
rect 352 338 368 358
rect 379 338 395 358
rect 407 304 423 358
rect 434 304 450 358
rect 462 212 478 358
rect 489 212 505 358
rect 520 158 536 358
rect 547 158 563 358
rect 574 158 590 358
rect 689 338 705 358
rect 716 338 732 358
rect 744 304 760 358
rect 771 304 787 358
rect 799 212 815 358
rect 826 212 842 358
rect 857 158 873 358
rect 884 158 900 358
rect 911 158 927 358
rect 1026 338 1042 358
rect 1053 338 1069 358
rect 1081 304 1097 358
rect 1108 304 1124 358
rect 1136 212 1152 358
rect 1163 212 1179 358
rect 1194 158 1210 358
rect 1221 158 1237 358
rect 1248 158 1264 358
rect 1371 337 1387 367
rect 1398 337 1414 367
<< pdiffcontact >>
rect 519 610 536 688
rect 352 398 368 456
rect 379 398 395 456
rect 407 398 423 555
rect 434 398 450 555
rect 462 398 478 610
rect 489 398 505 610
rect 516 398 536 610
rect 547 398 563 688
rect 574 398 590 688
rect 601 398 617 688
rect 628 398 644 688
rect 856 610 873 688
rect 689 398 705 456
rect 716 398 732 456
rect 744 398 760 555
rect 771 398 787 555
rect 799 398 815 610
rect 826 398 842 610
rect 853 398 873 610
rect 884 398 900 688
rect 911 398 927 688
rect 938 398 954 688
rect 965 398 981 688
rect 1193 610 1210 688
rect 1026 398 1042 456
rect 1053 398 1069 456
rect 1081 398 1097 555
rect 1108 398 1124 555
rect 1136 398 1152 610
rect 1163 398 1179 610
rect 1190 398 1210 610
rect 1221 398 1237 688
rect 1248 398 1264 688
rect 1275 398 1291 688
rect 1302 398 1318 688
rect 1371 413 1387 461
rect 1398 413 1414 461
<< psubstratetap >>
rect 326 66 342 82
rect 354 66 370 82
rect 382 66 398 82
rect 410 66 426 82
rect 438 66 454 82
rect 466 66 482 82
rect 494 66 510 82
rect 522 66 538 82
rect 550 66 567 82
rect 579 66 595 82
rect 607 66 623 82
rect 635 66 651 82
rect 663 66 679 82
rect 691 66 707 82
rect 719 66 735 82
rect 747 66 763 82
rect 775 66 791 82
rect 803 66 819 82
rect 831 66 847 82
rect 859 66 875 82
rect 887 66 904 82
rect 916 66 932 82
rect 944 66 960 82
rect 972 66 988 82
rect 1000 66 1016 82
rect 1028 66 1044 82
rect 1056 66 1072 82
rect 1084 66 1100 82
rect 1112 66 1128 82
rect 1140 66 1156 82
rect 1168 66 1184 82
rect 1196 66 1212 82
rect 1224 66 1241 82
rect 1253 66 1269 82
rect 1281 66 1297 82
rect 1309 66 1325 82
rect 1337 66 1353 82
rect 1365 66 1381 82
rect 1393 66 1409 82
rect 1421 66 1437 82
<< nsubstratetap >>
rect 214 720 230 736
rect 242 720 258 736
rect 270 720 286 736
rect 298 720 314 736
rect 326 720 342 736
rect 354 720 370 736
rect 382 720 398 736
rect 410 720 426 736
rect 438 720 454 736
rect 466 720 482 736
rect 494 720 510 736
rect 522 720 538 736
rect 550 720 567 736
rect 579 720 595 736
rect 607 720 623 736
rect 635 720 651 736
rect 663 720 679 736
rect 691 720 707 736
rect 719 720 735 736
rect 747 720 763 736
rect 775 720 791 736
rect 803 720 819 736
rect 831 720 847 736
rect 859 720 875 736
rect 887 720 904 736
rect 916 720 932 736
rect 944 720 960 736
rect 972 720 988 736
rect 1000 720 1016 736
rect 1028 720 1044 736
rect 1056 720 1072 736
rect 1084 720 1100 736
rect 1112 720 1128 736
rect 1140 720 1156 736
rect 1168 720 1184 736
rect 1196 720 1212 736
rect 1224 720 1241 736
rect 1253 720 1269 736
rect 1281 720 1297 736
rect 1309 720 1325 736
rect 1337 720 1353 736
rect 1365 720 1381 736
rect 1393 720 1409 736
rect 1421 720 1437 736
<< metal1 >>
rect 236 772 1356 782
rect 1400 772 1464 782
rect 236 749 1464 759
rect 200 720 214 736
rect 230 720 242 736
rect 258 720 270 736
rect 286 720 298 736
rect 314 720 326 736
rect 342 720 354 736
rect 370 720 382 736
rect 398 720 410 736
rect 426 720 438 736
rect 454 720 466 736
rect 482 720 494 736
rect 510 720 522 736
rect 538 720 550 736
rect 567 720 579 736
rect 595 720 607 736
rect 623 720 635 736
rect 651 720 663 736
rect 679 720 691 736
rect 707 720 719 736
rect 735 720 747 736
rect 763 720 775 736
rect 791 720 803 736
rect 819 720 831 736
rect 847 720 859 736
rect 875 720 887 736
rect 904 720 916 736
rect 932 720 944 736
rect 960 720 972 736
rect 988 720 1000 736
rect 1016 720 1028 736
rect 1044 720 1056 736
rect 1072 720 1084 736
rect 1100 720 1112 736
rect 1128 720 1140 736
rect 1156 720 1168 736
rect 1184 720 1196 736
rect 1212 720 1224 736
rect 1241 720 1253 736
rect 1269 720 1281 736
rect 1297 720 1309 736
rect 1325 720 1337 736
rect 1353 720 1365 736
rect 1381 720 1393 736
rect 1409 720 1421 736
rect 1437 720 1464 736
rect 200 711 1464 720
rect 352 456 368 711
rect 407 555 423 711
rect 462 610 478 711
rect 516 688 536 711
rect 574 688 590 711
rect 628 688 644 711
rect 516 610 519 688
rect 689 456 705 711
rect 744 555 760 711
rect 799 610 815 711
rect 853 688 873 711
rect 911 688 927 711
rect 965 688 981 711
rect 853 610 856 688
rect 1026 456 1042 711
rect 1081 555 1097 711
rect 1136 610 1152 711
rect 1190 688 1210 711
rect 1248 688 1264 711
rect 1302 688 1318 711
rect 1190 610 1193 688
rect 1380 522 1394 528
rect 1404 461 1414 711
rect 284 371 359 381
rect 270 359 284 369
rect 385 381 395 398
rect 385 371 414 381
rect 385 358 395 371
rect 440 382 450 398
rect 440 372 469 382
rect 440 358 450 372
rect 495 382 505 398
rect 495 372 527 382
rect 495 358 505 372
rect 553 383 563 398
rect 607 385 617 398
rect 553 373 606 383
rect 553 358 563 373
rect 667 371 696 381
rect 722 381 732 398
rect 722 371 751 381
rect 722 358 732 371
rect 777 382 787 398
rect 777 372 806 382
rect 777 358 787 372
rect 832 382 842 398
rect 832 372 864 382
rect 832 358 842 372
rect 890 383 900 398
rect 944 385 954 398
rect 890 373 944 383
rect 890 358 900 373
rect 1022 371 1033 381
rect 1059 381 1069 398
rect 1059 371 1088 381
rect 1059 358 1069 371
rect 1114 382 1124 398
rect 1114 372 1143 382
rect 1114 358 1124 372
rect 1169 382 1179 398
rect 1169 372 1201 382
rect 1169 358 1179 372
rect 1227 383 1237 398
rect 1281 385 1291 398
rect 1227 373 1279 383
rect 1227 358 1237 373
rect 1371 367 1381 413
rect 352 91 368 338
rect 407 91 423 304
rect 462 91 478 212
rect 520 91 536 158
rect 574 91 590 158
rect 689 91 705 338
rect 744 91 760 304
rect 799 91 815 212
rect 857 91 873 158
rect 911 91 927 158
rect 1026 91 1042 338
rect 1081 91 1097 304
rect 1136 91 1152 212
rect 1194 91 1210 158
rect 1248 91 1264 158
rect 1398 91 1408 337
rect 320 82 1464 91
rect 320 66 326 82
rect 342 66 354 82
rect 370 66 382 82
rect 398 66 410 82
rect 426 66 438 82
rect 454 66 466 82
rect 482 66 494 82
rect 510 66 522 82
rect 538 66 550 82
rect 567 66 579 82
rect 595 66 607 82
rect 623 66 635 82
rect 651 66 663 82
rect 679 66 691 82
rect 707 66 719 82
rect 735 66 747 82
rect 763 66 775 82
rect 791 66 803 82
rect 819 66 831 82
rect 847 66 859 82
rect 875 66 887 82
rect 904 66 916 82
rect 932 66 944 82
rect 960 66 972 82
rect 988 66 1000 82
rect 1016 66 1028 82
rect 1044 66 1056 82
rect 1072 66 1084 82
rect 1100 66 1112 82
rect 1128 66 1140 82
rect 1156 66 1168 82
rect 1184 66 1196 82
rect 1212 66 1224 82
rect 1241 66 1253 82
rect 1269 66 1281 82
rect 1297 66 1309 82
rect 1325 66 1337 82
rect 1353 66 1365 82
rect 1381 66 1393 82
rect 1409 66 1421 82
rect 1437 66 1464 82
rect 246 33 260 43
rect 620 43 1464 53
rect 260 20 653 30
rect 959 20 1464 30
rect 308 -3 1009 7
rect 1294 -3 1304 7
rect 1318 -3 1464 7
<< m2contact >>
rect 222 770 236 784
rect 1356 771 1370 785
rect 1386 771 1400 785
rect 222 746 236 760
rect 0 711 200 736
rect 1380 528 1394 542
rect 1357 447 1371 461
rect 270 369 284 383
rect 270 345 284 359
rect 606 371 620 385
rect 653 369 667 383
rect 944 371 958 385
rect 1008 369 1022 383
rect 1279 371 1293 385
rect 246 43 260 57
rect 606 41 620 55
rect 246 19 260 33
rect 653 18 667 32
rect 945 19 959 33
rect 246 -5 260 9
rect 270 -5 284 9
rect 294 -5 308 9
rect 1009 -5 1023 9
rect 1280 -5 1294 9
rect 1304 -5 1318 9
<< metal2 >>
rect 0 736 200 789
rect 223 784 235 789
rect 0 -10 200 711
rect 223 -10 235 746
rect 247 57 259 789
rect 271 383 283 789
rect 271 359 283 369
rect 247 33 259 43
rect 247 9 259 19
rect 271 9 283 345
rect 295 9 307 789
rect 1358 461 1370 771
rect 1386 542 1398 771
rect 1394 528 1398 542
rect 607 55 619 371
rect 654 32 666 369
rect 946 33 958 371
rect 1010 9 1022 369
rect 1281 9 1293 371
rect 1294 -5 1304 9
rect 247 -10 259 -5
rect 271 -10 283 -5
rect 295 -10 307 -5
<< labels >>
rlabel metal2 0 789 200 789 5 Vdd!
rlabel metal2 247 789 259 789 5 Test
rlabel metal2 271 789 283 789 5 Clock
rlabel metal2 295 789 307 789 5 nReset
rlabel metal2 247 -10 259 -10 1 Test
rlabel metal2 271 -10 283 -10 1 Clock
rlabel metal2 0 -10 200 -10 1 Vdd!
rlabel metal2 295 -10 307 -10 1 nReset
rlabel metal2 223 -10 235 -10 1 SDI
rlabel metal1 1464 711 1464 736 7 Vdd!
rlabel metal1 1464 749 1464 759 7 SDI
rlabel metal1 1464 772 1464 782 7 nSDO
rlabel metal1 1464 43 1464 53 7 ClockOut
rlabel metal1 1464 20 1464 30 7 TestOut
rlabel metal1 1464 -3 1464 7 7 nResetOut
rlabel metal1 1464 66 1464 91 7 GND!
<< end >>
