magic
tech c035u
timestamp 1386006835
use ../leftbuf/leftbuf leftbuf_0
timestamp 1386006472
transform 1 0 0 0 1 0
box 0 0 1464 799
use ../and2/and2 and2_0
timestamp 1385636468
transform 1 0 1464 0 1 0
box 0 0 120 799
use ../nand2/nand2 nand2_0
timestamp 1385998521
transform 1 0 1584 0 1 0
box 0 0 96 799
use ../nand3/nand3 nand3_0
timestamp 1385998574
transform 1 0 1680 0 1 0
box 0 0 120 799
use ../nand4/nand4 nand4_0
timestamp 1385998349
transform 1 0 1800 0 1 0
box 0 0 144 799
use ../nor2/nor2 nor2_0
timestamp 1385632928
transform 1 0 1944 0 1 0
box 0 0 120 799
use ../nor3/nor3 nor3_0
timestamp 1385633286
transform 1 0 2064 0 1 0
box 0 0 144 799
use ../or2/or2 or2_0
timestamp 1385633707
transform 1 0 2208 0 1 0
box 0 0 144 799
use ../mux2/mux2 mux2_0
timestamp 1385925694
transform 1 0 2352 0 1 0
box 0 0 192 799
use ../smux2/smux2 smux2_0
timestamp 1385926013
transform 1 0 2544 0 1 0
box 0 0 192 799
use ../smux3/smux3 smux3_0
timestamp 1385926127
transform 1 0 2736 0 1 0
box 0 0 288 799
use ../buffer/buffer buffer_0
timestamp 1385998845
transform 1 0 3024 0 1 0
box 0 0 120 799
use ../inv/inv inv_0
timestamp 1385924870
transform 1 0 3144 0 1 0
box 0 0 120 799
use ../trisbuf/trisbuf trisbuf_0
timestamp 1385926402
transform 1 0 3264 0 1 0
box 0 0 192 799
use ../rdtype/rdtype rdtype_0
timestamp 1386002196
transform 1 0 3456 0 1 0
box 0 0 432 799
use ../fulladder/fulladder fulladder_0
timestamp 1386001875
transform 1 0 3888 0 1 0
box 0 0 360 799
use ../halfadder/halfadder halfadder_0
timestamp 1385925245
transform 1 0 4248 0 1 0
box 0 0 312 799
use ../xor2/xor2 xor2_0
timestamp 1385932968
transform 1 0 4560 0 1 0
box 0 0 192 799
use ../tielow/tielow tielow_0
timestamp 1385999837
transform 1 0 4752 0 1 0
box 0 0 48 799
use ../tiehigh/tiehigh tiehigh_0
timestamp 1386006554
transform 1 0 4800 0 1 0
box 0 0 48 799
use ../rowcrosser/rowcrosser rowcrosser_0
timestamp 1386006577
transform 1 0 4848 0 1 0
box 0 0 48 799
use ../scandtype/scandtype scandtype_0
timestamp 1385994490
transform 1 0 4896 0 1 0
box 0 0 648 799
use ../scanreg/scanreg scanreg_0
timestamp 1386006598
transform 1 0 5544 0 1 0
box 0 0 768 799
use ../rightend/rightend rightend_0
timestamp 1386006533
transform 1 0 6312 0 1 0
box 0 0 320 799
<< end >>
