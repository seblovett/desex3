magic
tech c035u
timestamp 1386236433
<< nwell >>
rect 0 401 624 799
<< pwell >>
rect 0 0 624 401
<< polysilicon >>
rect 29 691 36 699
rect 59 691 66 699
rect 88 691 95 699
rect 115 691 122 699
rect 146 691 153 699
rect 259 691 266 719
rect 289 691 296 719
rect 340 704 407 711
rect 29 612 36 643
rect 59 599 66 643
rect 29 347 36 564
rect 59 347 66 583
rect 88 573 95 643
rect 115 591 122 643
rect 146 633 153 643
rect 149 617 153 633
rect 115 575 116 591
rect 88 347 95 557
rect 115 347 122 575
rect 146 393 153 617
rect 226 610 233 621
rect 148 377 153 393
rect 226 388 233 562
rect 259 486 266 643
rect 289 612 296 643
rect 342 612 349 623
rect 383 612 390 645
rect 400 624 407 704
rect 445 691 452 719
rect 503 691 510 719
rect 445 624 452 643
rect 400 617 452 624
rect 445 612 452 617
rect 289 486 296 564
rect 342 486 349 564
rect 383 486 390 564
rect 445 486 452 564
rect 503 532 510 643
rect 571 612 578 675
rect 29 282 36 317
rect 59 278 66 317
rect 88 309 95 317
rect 115 309 122 317
rect 146 282 153 377
rect 29 242 36 252
rect 146 244 153 252
rect 29 226 37 242
rect 226 225 233 372
rect 259 331 266 438
rect 289 402 296 438
rect 342 428 349 438
rect 358 412 370 419
rect 289 395 330 402
rect 323 358 330 395
rect 363 358 370 412
rect 383 410 390 438
rect 445 428 452 438
rect 383 403 411 410
rect 404 358 411 403
rect 445 358 452 412
rect 259 288 266 315
rect 323 288 330 328
rect 226 187 233 195
rect 259 161 266 258
rect 323 225 330 258
rect 363 225 370 328
rect 404 225 411 328
rect 445 255 452 328
rect 445 248 459 255
rect 445 225 459 232
rect 445 220 452 225
rect 503 220 510 516
rect 535 486 542 539
rect 535 358 542 438
rect 535 288 542 328
rect 259 110 266 131
rect 323 127 330 195
rect 363 128 370 195
rect 404 161 411 195
rect 445 161 452 190
rect 503 180 510 190
rect 503 142 510 150
rect 535 142 542 258
rect 571 227 578 564
rect 561 220 578 227
rect 568 190 575 195
rect 561 188 575 190
rect 568 180 575 188
rect 568 142 575 150
rect 404 120 411 131
rect 445 120 452 131
<< ndiffusion >>
rect 27 317 29 347
rect 36 317 38 347
rect 54 317 59 347
rect 66 317 88 347
rect 95 317 97 347
rect 113 317 115 347
rect 122 317 124 347
rect 27 252 29 282
rect 36 252 38 282
rect 144 252 146 282
rect 153 252 155 282
rect 318 328 323 358
rect 330 328 363 358
rect 370 328 377 358
rect 393 328 404 358
rect 411 328 445 358
rect 452 328 457 358
rect 254 258 259 288
rect 266 258 323 288
rect 330 258 341 288
rect 224 195 226 225
rect 233 195 238 225
rect 321 195 323 225
rect 330 195 363 225
rect 370 195 373 225
rect 533 258 535 288
rect 542 258 548 288
rect 254 131 259 161
rect 266 131 271 161
rect 437 190 445 220
rect 452 190 503 220
rect 510 190 514 220
rect 402 131 404 161
rect 411 131 445 161
rect 452 131 456 161
rect 565 150 568 180
rect 575 150 578 180
<< pdiffusion >>
rect 27 643 29 691
rect 36 643 38 691
rect 54 643 59 691
rect 66 643 68 691
rect 84 643 88 691
rect 95 643 97 691
rect 113 643 115 691
rect 122 643 125 691
rect 141 643 146 691
rect 153 643 156 691
rect 257 643 259 691
rect 266 643 268 691
rect 284 643 289 691
rect 296 643 298 691
rect 27 564 29 612
rect 36 564 38 612
rect 223 562 226 610
rect 233 562 238 610
rect 428 643 445 691
rect 452 643 462 691
rect 478 643 503 691
rect 510 643 513 691
rect 287 564 289 612
rect 296 564 324 612
rect 340 564 342 612
rect 349 564 359 612
rect 375 564 383 612
rect 390 564 392 612
rect 408 564 445 612
rect 452 564 454 612
rect 568 564 571 612
rect 578 564 588 612
rect 257 438 259 486
rect 266 438 269 486
rect 285 438 289 486
rect 296 438 298 486
rect 318 438 342 486
rect 349 438 357 486
rect 375 438 383 486
rect 390 438 392 486
rect 408 438 445 486
rect 452 438 455 486
rect 532 438 535 486
rect 542 438 548 486
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 202 86
rect 0 76 202 79
rect 218 76 230 86
rect 246 76 258 86
rect 274 76 286 86
rect 302 76 314 86
rect 330 76 342 86
rect 358 76 370 86
rect 386 76 398 86
rect 414 76 426 86
rect 443 76 455 86
rect 471 76 483 86
rect 499 76 511 86
rect 527 76 539 86
rect 556 76 568 86
rect 585 76 597 86
rect 614 76 624 86
<< nohmic >>
rect 0 743 202 746
rect 0 736 8 743
rect 24 736 36 743
rect 52 736 64 743
rect 80 736 92 743
rect 108 736 120 743
rect 136 736 148 743
rect 164 736 202 743
rect 218 736 230 746
rect 246 736 258 746
rect 274 736 286 746
rect 302 736 314 746
rect 330 736 342 746
rect 358 736 370 746
rect 386 736 398 746
rect 414 736 426 746
rect 442 736 454 746
rect 470 736 482 746
rect 498 736 510 746
rect 526 736 538 746
rect 554 736 566 746
rect 582 736 594 746
rect 610 736 624 746
<< ntransistor >>
rect 29 317 36 347
rect 59 317 66 347
rect 88 317 95 347
rect 115 317 122 347
rect 29 252 36 282
rect 146 252 153 282
rect 323 328 330 358
rect 363 328 370 358
rect 404 328 411 358
rect 445 328 452 358
rect 259 258 266 288
rect 323 258 330 288
rect 226 195 233 225
rect 323 195 330 225
rect 363 195 370 225
rect 535 258 542 288
rect 259 131 266 161
rect 445 190 452 220
rect 503 190 510 220
rect 404 131 411 161
rect 445 131 452 161
rect 568 150 575 180
<< ptransistor >>
rect 29 643 36 691
rect 59 643 66 691
rect 88 643 95 691
rect 115 643 122 691
rect 146 643 153 691
rect 259 643 266 691
rect 289 643 296 691
rect 29 564 36 612
rect 226 562 233 610
rect 445 643 452 691
rect 503 643 510 691
rect 289 564 296 612
rect 342 564 349 612
rect 383 564 390 612
rect 445 564 452 612
rect 571 564 578 612
rect 259 438 266 486
rect 289 438 296 486
rect 342 438 349 486
rect 383 438 390 486
rect 445 438 452 486
rect 535 438 542 486
<< polycontact >>
rect 324 695 340 711
rect 374 645 390 661
rect 59 583 75 599
rect 133 617 149 633
rect 116 575 132 591
rect 84 557 100 573
rect 132 377 148 393
rect 562 675 578 691
rect 526 539 542 555
rect 498 516 514 532
rect 217 372 233 388
rect 59 262 75 278
rect 37 226 53 242
rect 342 412 358 428
rect 445 412 461 428
rect 255 315 271 331
rect 447 232 463 248
rect 395 195 411 225
rect 526 328 542 358
rect 503 150 519 180
rect 552 190 568 220
rect 318 111 334 127
rect 359 111 376 128
<< ndiffcontact >>
rect 11 317 27 347
rect 38 317 54 347
rect 97 317 113 347
rect 124 317 140 347
rect 11 252 27 282
rect 38 252 54 282
rect 128 252 144 282
rect 155 252 175 282
rect 302 328 318 358
rect 377 328 393 358
rect 457 328 473 358
rect 238 258 254 288
rect 341 258 357 288
rect 208 195 224 225
rect 238 195 254 225
rect 305 195 321 225
rect 373 195 389 225
rect 517 258 533 288
rect 548 258 564 288
rect 238 131 254 161
rect 271 131 287 161
rect 421 190 437 220
rect 514 190 530 220
rect 386 131 402 161
rect 456 131 472 161
rect 549 150 565 180
rect 578 150 594 180
<< pdiffcontact >>
rect 11 643 27 691
rect 38 643 54 691
rect 68 643 84 691
rect 97 643 113 691
rect 125 643 141 691
rect 156 643 176 691
rect 241 643 257 691
rect 268 643 284 691
rect 298 643 314 691
rect 11 564 27 612
rect 38 564 54 612
rect 207 562 223 610
rect 238 562 254 610
rect 412 643 428 691
rect 462 643 478 691
rect 513 643 529 691
rect 271 564 287 612
rect 324 564 340 612
rect 359 564 375 612
rect 392 564 408 612
rect 454 564 470 612
rect 552 564 568 612
rect 588 564 604 612
rect 241 438 257 486
rect 269 438 285 486
rect 298 438 318 486
rect 357 438 375 486
rect 392 438 408 486
rect 455 438 471 486
rect 516 438 532 486
rect 548 438 565 486
<< psubstratetap >>
rect 128 216 144 232
rect 208 166 224 182
rect 6 79 22 95
rect 34 79 50 95
rect 62 79 78 95
rect 90 79 106 95
rect 118 79 134 95
rect 146 79 162 95
rect 202 76 218 92
rect 230 76 246 92
rect 258 76 274 92
rect 286 76 302 92
rect 314 76 330 92
rect 342 76 358 92
rect 370 76 386 92
rect 398 76 414 92
rect 426 76 443 92
rect 455 76 471 92
rect 483 76 499 92
rect 511 76 527 92
rect 539 76 556 92
rect 568 76 585 92
rect 597 76 614 92
<< nsubstratetap >>
rect 8 727 24 743
rect 36 727 52 743
rect 64 727 80 743
rect 92 727 108 743
rect 120 727 136 743
rect 148 727 164 743
rect 202 730 218 746
rect 230 730 246 746
rect 258 730 274 746
rect 286 730 302 746
rect 314 730 330 746
rect 342 730 358 746
rect 370 730 386 746
rect 398 730 414 746
rect 426 730 442 746
rect 454 730 470 746
rect 482 730 498 746
rect 510 730 526 746
rect 538 730 554 746
rect 566 730 582 746
rect 594 730 610 746
<< metal1 >>
rect 0 782 624 792
rect 0 759 118 769
rect 192 759 506 769
rect 522 759 624 769
rect 0 743 202 746
rect 0 727 8 743
rect 24 727 36 743
rect 52 727 64 743
rect 80 727 92 743
rect 108 727 120 743
rect 136 727 148 743
rect 164 730 202 743
rect 218 730 230 746
rect 246 730 258 746
rect 274 730 286 746
rect 302 730 314 746
rect 330 730 342 746
rect 358 730 370 746
rect 386 730 398 746
rect 414 730 426 746
rect 442 730 454 746
rect 470 730 482 746
rect 498 730 510 746
rect 526 730 538 746
rect 554 730 566 746
rect 582 730 594 746
rect 610 730 624 746
rect 164 727 624 730
rect 0 721 624 727
rect 11 691 27 721
rect 41 701 110 711
rect 41 691 51 701
rect 100 691 110 701
rect 125 691 141 721
rect 11 612 27 643
rect 71 629 81 643
rect 71 619 133 629
rect 54 583 59 599
rect 41 380 132 390
rect 41 347 51 380
rect 159 385 169 643
rect 207 634 223 721
rect 241 691 257 721
rect 268 701 324 711
rect 268 691 284 701
rect 462 701 562 711
rect 462 691 478 701
rect 562 691 578 695
rect 207 633 224 634
rect 298 633 314 643
rect 207 621 314 633
rect 324 645 374 655
rect 207 610 223 621
rect 271 612 287 621
rect 207 511 223 562
rect 324 612 340 645
rect 412 633 428 643
rect 513 633 529 643
rect 588 633 604 721
rect 359 623 604 633
rect 359 612 375 623
rect 454 612 470 623
rect 588 612 604 623
rect 238 549 254 562
rect 324 549 340 564
rect 238 539 340 549
rect 392 554 408 564
rect 392 544 526 554
rect 298 516 458 526
rect 474 516 498 526
rect 552 526 568 564
rect 514 516 568 526
rect 207 501 285 511
rect 269 486 285 501
rect 298 486 318 516
rect 588 506 604 564
rect 357 496 471 506
rect 357 486 375 496
rect 455 486 471 496
rect 516 496 604 506
rect 516 486 532 496
rect 471 438 516 486
rect 241 428 257 438
rect 392 428 408 438
rect 548 428 565 438
rect 241 418 342 428
rect 358 418 408 428
rect 461 418 565 428
rect 256 390 393 402
rect 159 375 217 385
rect 73 357 137 367
rect 14 307 24 317
rect 73 307 83 357
rect 127 347 137 357
rect 14 297 83 307
rect 54 262 59 278
rect 11 101 27 252
rect 97 101 113 317
rect 159 282 169 375
rect 256 353 269 390
rect 377 358 393 390
rect 208 341 269 353
rect 208 288 224 341
rect 255 314 271 315
rect 473 328 526 358
rect 302 318 318 328
rect 302 308 594 318
rect 208 258 238 288
rect 357 278 517 288
rect 128 232 144 252
rect 128 101 144 216
rect 208 225 224 258
rect 238 247 254 258
rect 548 248 564 258
rect 238 235 437 247
rect 254 195 305 225
rect 389 195 395 225
rect 421 220 437 235
rect 463 232 564 248
rect 208 182 224 195
rect 530 190 552 220
rect 578 180 594 308
rect 208 161 224 166
rect 208 131 238 161
rect 287 151 386 161
rect 519 150 549 180
rect 208 101 226 131
rect 317 111 318 127
rect 456 121 472 131
rect 376 111 472 121
rect 0 95 624 101
rect 0 79 6 95
rect 22 79 34 95
rect 50 79 62 95
rect 78 79 90 95
rect 106 79 118 95
rect 134 79 146 95
rect 162 92 624 95
rect 162 79 202 92
rect 0 76 202 79
rect 218 76 230 92
rect 246 76 258 92
rect 274 76 286 92
rect 302 76 314 92
rect 330 76 342 92
rect 358 76 370 92
rect 386 76 398 92
rect 414 76 426 92
rect 443 76 455 92
rect 471 76 483 92
rect 499 76 511 92
rect 527 76 539 92
rect 556 76 568 92
rect 585 76 597 92
rect 614 76 624 92
rect 0 53 255 63
rect 271 53 624 63
rect 0 30 39 40
rect 53 30 624 40
rect 0 7 301 17
rect 317 7 624 17
<< m2contact >>
rect 118 757 132 771
rect 506 756 522 772
rect 118 591 132 605
rect 85 543 99 557
rect 562 695 578 711
rect 458 516 474 532
rect 39 212 53 226
rect 255 298 271 314
rect 301 111 317 127
rect 255 50 271 66
rect 39 28 53 42
rect 301 4 317 20
<< metal2 >>
rect 96 557 108 799
rect 119 605 131 757
rect 99 543 108 557
rect 40 42 52 212
rect 96 0 108 543
rect 460 532 472 799
rect 508 772 520 799
rect 508 711 520 756
rect 508 695 562 711
rect 255 66 271 298
rect 301 20 317 111
rect 460 0 472 516
rect 508 0 520 695
<< labels >>
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal2 96 799 108 799 5 D
rlabel metal1 0 76 0 101 1 GND!
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 3 Clock
rlabel metal2 96 0 108 0 1 D
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal2 460 799 472 799 5 nQ
rlabel metal2 460 0 472 0 1 nQ
rlabel metal2 508 799 520 799 5 Q
rlabel metal2 508 0 520 0 1 Q
rlabel metal1 624 782 624 792 7 ScanReturn
rlabel metal1 624 759 624 769 7 Q
rlabel metal1 624 76 624 101 7 GND!
rlabel metal1 624 53 624 63 7 Clock
rlabel metal1 624 30 624 40 7 Test
rlabel metal1 624 7 624 17 7 nReset
rlabel metal1 624 721 624 746 7 Vdd!
<< end >>
