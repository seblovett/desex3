magic
tech c035u
timestamp 1385581317
<< nwell >>
rect 0 460 188 659
<< polysilicon >>
rect 29 604 36 612
rect 59 604 66 612
rect 88 604 95 612
rect 115 604 122 612
rect 146 604 153 612
rect 29 525 36 556
rect 59 512 66 556
rect 29 270 36 477
rect 59 270 66 496
rect 88 486 95 556
rect 115 504 122 556
rect 146 546 153 556
rect 149 530 153 546
rect 115 488 116 504
rect 88 270 95 470
rect 115 270 122 488
rect 146 316 153 530
rect 148 300 153 316
rect 29 209 36 244
rect 59 205 66 244
rect 88 236 95 244
rect 115 236 122 244
rect 146 209 153 300
rect 29 173 36 183
rect 146 175 153 183
rect 29 157 37 173
<< ndiffusion >>
rect 27 244 29 270
rect 36 244 38 270
rect 54 244 59 270
rect 66 244 88 270
rect 95 244 97 270
rect 113 244 115 270
rect 122 244 124 270
rect 27 183 29 209
rect 36 183 38 209
rect 144 183 146 209
rect 153 183 155 209
<< pdiffusion >>
rect 27 556 29 604
rect 36 556 38 604
rect 54 556 59 604
rect 66 556 68 604
rect 84 556 88 604
rect 95 556 97 604
rect 113 556 115 604
rect 122 556 125 604
rect 141 556 146 604
rect 153 556 156 604
rect 27 477 29 525
rect 36 477 38 525
<< pohmic >>
rect 0 2 6 9
rect 22 2 34 9
rect 50 2 62 9
rect 78 2 90 9
rect 106 2 118 9
rect 134 2 146 9
rect 162 2 188 9
rect 0 -1 188 2
<< nohmic >>
rect 0 656 188 659
rect 0 649 8 656
rect 24 649 36 656
rect 52 649 64 656
rect 80 649 92 656
rect 108 649 120 656
rect 136 649 148 656
rect 164 649 188 656
<< ntransistor >>
rect 29 244 36 270
rect 59 244 66 270
rect 88 244 95 270
rect 115 244 122 270
rect 29 183 36 209
rect 146 183 153 209
<< ptransistor >>
rect 29 556 36 604
rect 59 556 66 604
rect 88 556 95 604
rect 115 556 122 604
rect 146 556 153 604
rect 29 477 36 525
<< polycontact >>
rect 59 496 75 512
rect 133 530 149 546
rect 116 488 132 504
rect 84 470 100 486
rect 132 300 148 316
rect 59 189 75 205
rect 37 157 53 173
<< ndiffcontact >>
rect 11 244 27 270
rect 38 244 54 270
rect 97 244 113 270
rect 124 244 140 270
rect 11 183 27 209
rect 38 183 54 209
rect 128 183 144 209
rect 155 183 171 209
<< pdiffcontact >>
rect 11 556 27 604
rect 38 556 54 604
rect 68 556 84 604
rect 97 556 113 604
rect 125 556 141 604
rect 156 556 172 604
rect 11 477 27 525
rect 38 477 54 525
<< psubstratetap >>
rect 6 2 22 18
rect 34 2 50 18
rect 62 2 78 18
rect 90 2 106 18
rect 118 2 134 18
rect 146 2 162 18
<< nsubstratetap >>
rect 8 640 24 656
rect 36 640 52 656
rect 64 640 80 656
rect 92 640 108 656
rect 120 640 136 656
rect 148 640 164 656
<< metal1 >>
rect 0 695 188 705
rect 0 672 118 682
rect 0 656 188 659
rect 0 640 8 656
rect 24 640 36 656
rect 52 640 64 656
rect 80 640 92 656
rect 108 640 120 656
rect 136 640 148 656
rect 164 640 188 656
rect 0 634 188 640
rect 11 604 27 634
rect 41 614 110 624
rect 41 604 51 614
rect 100 604 110 614
rect 125 604 141 634
rect 11 525 27 556
rect 71 542 81 556
rect 71 532 133 542
rect 54 496 59 512
rect 159 385 169 556
rect 159 375 188 385
rect 41 303 132 313
rect 41 270 51 303
rect 73 280 137 290
rect 14 234 24 244
rect 73 234 83 280
rect 127 270 137 280
rect 14 224 83 234
rect 54 189 59 205
rect 11 24 27 183
rect 97 24 113 244
rect 159 209 169 375
rect 128 24 144 183
rect 0 18 188 24
rect 0 2 6 18
rect 22 2 34 18
rect 50 2 62 18
rect 78 2 90 18
rect 106 2 118 18
rect 134 2 146 18
rect 162 2 188 18
rect 0 -1 188 2
rect 0 -24 188 -14
rect 0 -47 39 -37
rect 53 -47 188 -37
rect 0 -70 188 -60
<< m2contact >>
rect 118 670 132 684
rect 118 504 132 518
rect 85 456 99 470
rect 39 143 53 157
rect 39 -49 53 -35
<< metal2 >>
rect 96 470 108 709
rect 119 518 131 670
rect 99 456 108 470
rect 40 -35 52 143
rect 96 -74 108 456
<< labels >>
rlabel metal1 0 -1 0 24 1 GND!
rlabel metal1 0 -70 0 -60 2 nReset
rlabel metal1 0 -47 0 -37 3 Test
rlabel metal1 0 -24 0 -14 3 Clock
rlabel metal1 0 634 0 659 3 Vdd!
rlabel metal1 0 672 0 682 3 Scan
rlabel metal1 0 695 0 705 4 ScanReturn
rlabel metal1 188 -24 188 -14 7 Clock
rlabel metal1 188 -47 188 -37 7 Test
rlabel metal1 188 -70 188 -60 8 nReset
rlabel metal1 188 -1 188 24 7 GND!
rlabel metal2 96 -74 108 -74 1 D
rlabel metal2 96 709 108 709 5 D
rlabel metal1 188 375 188 385 7 M
rlabel metal1 188 634 188 659 7 Vdd!
rlabel metal1 188 695 188 705 6 ScanReturn
<< end >>
