magic
tech c035u
timestamp 1386237216
<< nwell >>
rect 0 401 216 799
<< pwell >>
rect 0 0 216 401
<< polysilicon >>
rect 142 627 149 636
rect 100 558 117 565
rect 67 548 74 556
rect 110 548 117 558
rect 67 490 74 500
rect 33 469 40 477
rect 110 478 117 500
rect 142 490 149 579
rect 33 391 40 421
rect 33 365 40 375
rect 33 327 40 335
rect 67 330 74 474
rect 67 304 74 314
rect 110 304 117 328
rect 67 266 74 274
rect 110 264 117 274
rect 142 238 149 474
rect 142 200 149 208
<< ndiffusion >>
rect 31 335 33 365
rect 40 335 42 365
rect 61 274 67 304
rect 74 274 110 304
rect 117 274 119 304
rect 123 208 124 238
rect 140 208 142 238
rect 149 208 151 238
<< pdiffusion >>
rect 140 579 142 627
rect 149 579 151 627
rect 63 500 67 548
rect 74 500 110 548
rect 117 500 119 548
rect 31 421 33 469
rect 40 421 42 469
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 174 86
rect 190 76 216 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
rect 50 736 62 746
rect 78 736 90 746
rect 106 736 118 746
rect 134 736 146 746
rect 162 736 174 746
rect 190 736 216 746
<< ntransistor >>
rect 33 335 40 365
rect 67 274 74 304
rect 110 274 117 304
rect 142 208 149 238
<< ptransistor >>
rect 142 579 149 627
rect 67 500 74 548
rect 110 500 117 548
rect 33 421 40 469
<< polycontact >>
rect 84 558 100 574
rect 57 474 74 490
rect 32 375 48 391
rect 58 314 74 330
rect 142 474 158 490
rect 110 248 126 264
<< ndiffcontact >>
rect 15 335 31 365
rect 42 335 58 365
rect 45 274 61 304
rect 119 274 135 304
rect 124 208 140 238
rect 151 208 167 238
<< pdiffcontact >>
rect 123 579 140 627
rect 151 579 168 627
rect 45 500 63 548
rect 119 500 135 548
rect 15 421 31 469
rect 42 421 58 469
<< psubstratetap >>
rect 15 300 31 316
rect 15 272 31 288
rect 15 244 31 260
rect 15 216 31 232
rect 15 188 31 204
rect 15 160 31 176
rect 15 132 31 148
rect 15 104 31 120
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
rect 174 76 190 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
rect 62 730 78 746
rect 90 730 106 746
rect 118 730 134 746
rect 146 730 162 746
rect 174 730 190 746
<< metal1 >>
rect 0 782 216 792
rect 0 759 216 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 62 746
rect 78 730 90 746
rect 106 730 118 746
rect 134 730 146 746
rect 162 730 174 746
rect 190 730 216 746
rect 0 721 216 730
rect 15 469 31 721
rect 45 720 88 721
rect 45 548 63 720
rect 151 627 168 721
rect 110 626 123 627
rect 84 579 123 626
rect 84 574 100 579
rect 42 474 57 490
rect 42 469 58 474
rect 15 316 31 335
rect 42 314 58 335
rect 15 288 31 300
rect 15 260 31 272
rect 15 232 31 244
rect 15 204 31 216
rect 15 176 31 188
rect 15 148 31 160
rect 15 120 31 132
rect 15 101 31 104
rect 45 101 61 274
rect 84 238 100 558
rect 119 434 132 500
rect 142 473 158 474
rect 119 417 168 434
rect 119 304 132 417
rect 126 248 127 264
rect 84 208 124 238
rect 151 101 167 208
rect 0 92 216 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 174 92
rect 190 76 216 92
rect 0 53 216 63
rect 0 30 216 40
rect 0 7 216 17
<< m2contact >>
rect 16 375 32 391
rect 142 457 158 473
rect 168 417 182 434
rect 127 248 143 264
<< metal2 >>
rect 24 391 36 799
rect 32 375 36 391
rect 24 0 36 375
rect 96 473 108 799
rect 96 457 142 473
rect 96 264 108 457
rect 168 434 180 799
rect 96 248 127 264
rect 96 0 108 248
rect 168 0 180 417
<< labels >>
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 76 0 101 3 GND!
rlabel metal2 24 0 36 0 1 A
rlabel metal2 24 799 36 799 5 A
rlabel metal2 96 799 108 799 5 Enable
rlabel metal2 96 0 108 0 1 Enable
rlabel metal2 168 0 180 0 1 Y
rlabel metal2 168 799 180 799 5 Y
rlabel metal1 216 7 216 17 8 nReset
rlabel metal1 216 30 216 40 7 Test
rlabel metal1 216 53 216 63 7 Clock
rlabel metal1 216 782 216 792 6 ScanReturn
rlabel metal1 216 759 216 769 7 Scan
rlabel metal1 216 721 216 746 7 Vdd!
rlabel metal1 216 76 216 101 7 GND!
<< end >>
