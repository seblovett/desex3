magic
tech c035u
timestamp 1385920833
<< nwell >>
rect 0 402 185 746
<< polysilicon >>
rect 30 630 37 638
rect 57 630 64 638
rect 88 630 95 638
rect 30 505 37 582
rect 57 549 64 582
rect 88 572 95 582
rect 150 581 159 588
rect 57 505 64 533
rect 30 406 37 457
rect 28 399 37 406
rect 28 397 35 399
rect 28 379 35 381
rect 28 372 37 379
rect 30 366 37 372
rect 57 366 64 457
rect 88 366 95 556
rect 122 505 129 513
rect 152 505 159 581
rect 122 447 129 457
rect 30 293 37 336
rect 57 293 64 336
rect 88 293 95 345
rect 122 335 129 431
rect 152 335 159 457
rect 122 297 129 305
rect 152 287 159 305
rect 148 280 159 287
rect 30 255 37 263
rect 57 255 64 263
rect 88 255 95 263
<< ndiffusion >>
rect 27 336 30 366
rect 37 336 57 366
rect 64 336 66 366
rect 120 305 122 335
rect 129 305 133 335
rect 149 305 152 335
rect 159 305 161 335
rect 27 263 30 293
rect 37 263 39 293
rect 55 263 57 293
rect 64 263 66 293
rect 82 263 88 293
rect 95 263 97 293
<< pdiffusion >>
rect 28 582 30 630
rect 37 582 39 630
rect 55 582 57 630
rect 64 582 66 630
rect 82 582 88 630
rect 95 582 97 630
rect 28 457 30 505
rect 37 457 57 505
rect 64 457 67 505
rect 119 457 122 505
rect 129 457 152 505
rect 159 457 161 505
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 185 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
rect 50 736 62 746
rect 78 736 90 746
rect 106 736 118 746
rect 134 736 146 746
rect 162 736 185 746
<< ntransistor >>
rect 30 336 37 366
rect 57 336 64 366
rect 122 305 129 335
rect 152 305 159 335
rect 30 263 37 293
rect 57 263 64 293
rect 88 263 95 293
<< ptransistor >>
rect 30 582 37 630
rect 57 582 64 630
rect 88 582 95 630
rect 30 457 37 505
rect 57 457 64 505
rect 122 457 129 505
rect 152 457 159 505
<< polycontact >>
rect 134 581 150 597
rect 80 556 96 572
rect 48 533 64 549
rect 19 381 35 397
rect 113 431 129 447
rect 88 345 104 366
rect 132 263 148 287
<< ndiffcontact >>
rect 11 336 27 366
rect 66 336 82 366
rect 104 305 120 335
rect 133 305 149 335
rect 161 305 177 335
rect 11 263 27 293
rect 39 263 55 293
rect 66 263 82 293
rect 97 263 113 293
<< pdiffcontact >>
rect 12 582 28 630
rect 39 582 55 630
rect 66 582 82 630
rect 97 582 113 630
rect 12 457 28 505
rect 67 457 83 505
rect 103 457 119 505
rect 161 457 177 505
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
rect 62 730 78 746
rect 90 730 106 746
rect 118 730 134 746
rect 146 730 162 746
<< metal1 >>
rect 0 782 185 792
rect 0 759 185 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 62 746
rect 78 730 90 746
rect 106 730 118 746
rect 134 730 146 746
rect 162 730 185 746
rect 0 721 185 730
rect 12 630 28 721
rect 66 630 82 721
rect 113 582 134 596
rect 12 505 28 582
rect 42 569 52 582
rect 42 559 80 569
rect 48 532 64 533
rect 161 505 178 721
rect 119 457 149 467
rect 177 457 178 505
rect 67 445 83 457
rect 45 433 113 445
rect 19 397 35 398
rect 11 293 27 336
rect 45 293 55 433
rect 139 394 149 457
rect 82 345 88 366
rect 139 335 149 378
rect 66 305 104 324
rect 66 293 82 305
rect 113 263 132 287
rect 11 101 27 263
rect 66 101 82 263
rect 161 101 177 305
rect 0 92 185 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 185 92
rect 0 53 185 63
rect 0 30 185 40
rect 0 7 185 17
<< m2contact >>
rect 48 516 64 532
rect 19 398 35 414
rect 133 378 149 394
<< metal2 >>
rect 19 414 31 799
rect 48 532 60 799
rect 19 0 31 398
rect 48 0 60 516
rect 137 394 149 799
rect 137 0 149 378
<< labels >>
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 0 76 0 101 3 GND!
rlabel metal2 137 0 149 0 1 Y
rlabel metal2 19 0 31 0 1 A
rlabel metal2 48 0 60 0 1 B
rlabel metal1 185 7 185 17 8 nReset
rlabel metal1 185 30 185 40 7 Test
rlabel metal1 185 53 185 63 7 Clock
rlabel metal1 185 76 185 101 7 GND!
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal2 19 799 31 799 5 A
rlabel metal2 48 799 60 799 5 B
rlabel metal2 137 799 149 799 5 Y
<< end >>
