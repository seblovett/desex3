magic
tech c035u
timestamp 1384736574
<< nwell >>
rect 18 310 392 610
rect 19 298 392 310
rect 19 240 393 298
<< polysilicon >>
rect 37 436 44 506
rect 71 496 78 543
rect 124 496 131 579
rect 204 501 260 508
rect 204 496 211 501
rect 253 496 260 501
rect 294 496 301 610
rect 367 496 374 610
rect 37 102 44 388
rect 71 352 78 448
rect 124 436 131 448
rect 163 436 170 444
rect 204 436 211 446
rect 253 436 260 448
rect 124 352 131 388
rect 163 352 170 388
rect 204 352 211 388
rect 253 352 260 388
rect 294 378 301 448
rect 367 436 374 480
rect 71 150 78 304
rect 124 198 131 304
rect 163 294 170 304
rect 163 198 170 278
rect 204 198 211 304
rect 253 294 260 304
rect 253 198 260 278
rect 124 150 131 169
rect 37 23 44 72
rect 71 60 78 120
rect 124 102 131 120
rect 163 102 170 169
rect 204 102 211 169
rect 253 131 260 169
rect 253 102 260 115
rect 294 102 301 362
rect 326 352 333 388
rect 326 198 333 304
rect 326 152 333 182
rect 71 22 78 30
rect 124 23 131 72
rect 163 40 170 72
rect 204 60 211 72
rect 253 60 260 72
rect 294 61 301 72
rect 204 22 211 30
rect 253 22 260 30
rect 294 23 301 31
rect 326 23 333 122
rect 367 102 374 388
rect 367 61 374 72
rect 367 23 374 31
<< ndiffusion >>
rect 99 169 124 198
rect 131 169 163 198
rect 170 182 177 198
rect 193 182 204 198
rect 170 169 204 182
rect 211 169 253 198
rect 260 182 265 198
rect 260 169 281 182
rect 66 120 71 150
rect 78 120 124 150
rect 131 134 142 150
rect 131 120 158 134
rect 35 72 37 102
rect 44 72 50 102
rect 324 136 326 152
rect 308 122 326 136
rect 333 129 344 152
rect 333 122 360 129
rect 119 72 124 102
rect 131 72 163 102
rect 170 72 173 102
rect 243 72 253 102
rect 260 72 294 102
rect 301 72 305 102
rect 66 30 71 60
rect 78 44 103 60
rect 78 30 119 44
rect 202 44 204 60
rect 186 30 204 44
rect 211 30 253 60
rect 260 30 264 60
rect 361 31 367 61
rect 374 31 384 61
<< pdiffusion >>
rect 65 448 71 496
rect 78 448 102 496
rect 118 448 124 496
rect 131 470 149 496
rect 131 448 133 470
rect 34 388 37 436
rect 44 409 62 436
rect 44 388 46 409
rect 250 448 253 496
rect 260 448 270 496
rect 286 448 294 496
rect 301 470 320 496
rect 301 448 304 470
rect 121 419 124 436
rect 105 388 124 419
rect 131 409 163 436
rect 131 388 135 409
rect 151 388 163 409
rect 170 388 183 436
rect 201 388 204 436
rect 211 404 253 436
rect 211 388 234 404
rect 250 388 253 404
rect 260 419 262 436
rect 260 388 273 419
rect 348 405 367 436
rect 364 388 367 405
rect 374 388 376 436
rect 49 326 71 352
rect 65 304 71 326
rect 78 304 105 352
rect 121 304 124 352
rect 131 304 134 352
rect 150 304 163 352
rect 170 304 183 352
rect 201 304 204 352
rect 211 326 253 352
rect 211 304 226 326
rect 242 304 253 326
rect 260 304 263 352
rect 323 304 326 352
rect 333 326 351 352
rect 333 304 335 326
<< ntransistor >>
rect 124 169 131 198
rect 163 169 170 198
rect 204 169 211 198
rect 253 169 260 198
rect 71 120 78 150
rect 124 120 131 150
rect 37 72 44 102
rect 326 122 333 152
rect 124 72 131 102
rect 163 72 170 102
rect 253 72 260 102
rect 294 72 301 102
rect 71 30 78 60
rect 204 30 211 60
rect 253 30 260 60
rect 367 31 374 61
<< ptransistor >>
rect 71 448 78 496
rect 124 448 131 496
rect 37 388 44 436
rect 253 448 260 496
rect 294 448 301 496
rect 124 388 131 436
rect 163 388 170 436
rect 204 388 211 436
rect 253 388 260 436
rect 367 388 374 436
rect 71 304 78 352
rect 124 304 131 352
rect 163 304 170 352
rect 204 304 211 352
rect 253 304 260 352
rect 326 304 333 352
<< polycontact >>
rect 116 579 141 604
rect 62 543 105 568
rect 29 506 54 531
rect 195 480 211 496
rect 195 446 211 462
rect 358 480 374 496
rect 317 388 333 404
rect 289 362 305 378
rect 158 278 174 294
rect 253 278 269 294
rect 253 115 269 131
rect 317 182 333 198
rect 195 72 211 102
rect 159 23 176 40
rect 294 31 310 61
rect 358 72 374 102
<< ndiffcontact >>
rect 83 169 99 198
rect 177 182 193 220
rect 265 182 281 198
rect 50 120 66 150
rect 142 134 158 150
rect 19 72 35 102
rect 50 72 66 102
rect 308 136 324 152
rect 344 129 360 152
rect 103 72 119 102
rect 173 72 189 102
rect 227 72 243 102
rect 305 72 321 102
rect 50 30 66 60
rect 103 44 119 60
rect 186 44 202 60
rect 264 30 280 60
rect 345 31 361 61
rect 384 31 400 61
<< pdiffcontact >>
rect 49 448 65 496
rect 102 448 118 496
rect 133 448 149 470
rect 18 388 34 436
rect 46 388 62 409
rect 234 448 250 496
rect 270 448 286 496
rect 304 448 320 470
rect 105 419 121 436
rect 135 388 151 409
rect 183 388 201 436
rect 234 388 250 404
rect 262 419 278 436
rect 348 388 364 405
rect 376 388 392 436
rect 49 304 65 326
rect 105 304 121 352
rect 134 304 150 352
rect 183 304 201 352
rect 226 304 242 326
rect 263 304 279 352
rect 307 304 323 352
rect 335 304 351 326
<< psubstratetap >>
rect 136 212 154 228
<< nsubstratetap >>
rect 137 249 155 265
<< metal1 >>
rect 0 579 116 604
rect 141 579 406 604
rect 0 543 62 568
rect 105 543 406 568
rect 0 506 29 531
rect 54 506 406 531
rect 118 480 195 496
rect 49 436 65 448
rect 133 436 149 448
rect 34 419 105 436
rect 121 419 149 436
rect 159 446 195 462
rect 286 480 358 496
rect 159 409 172 446
rect 234 436 250 448
rect 304 436 320 448
rect 62 388 135 409
rect 151 388 172 409
rect 201 419 262 436
rect 278 419 376 436
rect 250 388 317 404
rect 18 352 34 388
rect 348 378 364 388
rect 134 362 289 378
rect 305 362 364 378
rect 134 352 150 362
rect 376 352 392 388
rect 18 336 105 352
rect 18 310 34 336
rect 19 268 34 310
rect 201 336 263 352
rect 279 336 307 352
rect 323 336 392 352
rect 49 294 65 304
rect 226 294 242 304
rect 335 294 351 304
rect 49 278 158 294
rect 174 278 242 294
rect 269 278 351 294
rect 376 268 392 336
rect 0 265 407 268
rect 0 249 137 265
rect 155 249 407 265
rect 0 243 407 249
rect 0 228 407 233
rect 0 212 136 228
rect 154 220 407 228
rect 154 212 177 220
rect 0 208 177 212
rect 19 150 35 208
rect 193 208 407 220
rect 281 182 317 198
rect 99 169 400 172
rect 83 162 400 169
rect 142 150 308 152
rect 19 120 50 150
rect 158 141 308 150
rect 66 120 243 122
rect 19 112 243 120
rect 344 126 360 129
rect 269 115 360 126
rect 19 102 35 112
rect 227 102 243 112
rect 66 72 103 102
rect 189 72 195 102
rect 321 72 358 102
rect 19 60 35 72
rect 384 61 400 162
rect 19 30 50 60
rect 119 50 186 60
rect 176 30 264 34
rect 310 31 345 61
rect 176 23 280 30
<< labels >>
rlabel metal1 0 243 0 268 3 Vdd!
rlabel metal1 0 208 0 233 3 GND!
rlabel metal1 0 579 0 604 3 nRst
rlabel metal1 0 543 0 568 3 Clk
rlabel metal1 0 506 0 531 3 D
rlabel metal1 407 243 407 268 7 Vdd!
rlabel metal1 407 208 407 233 7 GND!
rlabel metal1 406 579 406 604 7 nRst
rlabel metal1 406 543 406 568 7 Clk
rlabel metal1 406 506 406 531 7 D
rlabel polysilicon 367 610 374 610 5 Q
rlabel polysilicon 294 610 301 610 5 nQ
<< end >>
