magic
tech c035u
timestamp 1386341366
<< metal1 >>
rect 205 836 286 846
rect 85 810 261 820
rect 325 810 359 820
rect 373 810 479 820
<< m2contact >>
rect 191 833 205 847
rect 286 834 300 848
rect 71 807 85 821
rect 261 808 275 822
rect 311 808 325 822
rect 359 808 373 822
rect 479 808 493 822
<< metal2 >>
rect 24 799 36 862
rect 72 799 84 807
rect 144 799 156 862
rect 192 799 204 833
rect 264 822 276 862
rect 288 848 300 862
rect 275 808 276 822
rect 264 799 276 808
rect 288 799 300 834
rect 312 822 324 862
rect 312 799 324 808
rect 360 799 372 808
rect 408 799 420 862
rect 480 799 492 808
rect 528 799 540 862
use inv inv_0
timestamp 1386238110
transform 1 0 0 0 1 0
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 120 0 1 0
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 240 0 1 0
box 0 0 96 799
use inv inv_2
timestamp 1386238110
transform 1 0 336 0 1 0
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 456 0 1 0
box 0 0 120 799
<< labels >>
rlabel metal2 24 862 36 862 5 NA
rlabel metal2 144 862 156 862 5 NB
rlabel metal2 264 862 276 862 5 A
rlabel metal2 288 862 300 862 5 B
rlabel metal2 312 862 324 862 5 Y
rlabel metal2 408 862 420 862 5 n1
rlabel metal2 528 862 540 862 5 n2
<< end >>
