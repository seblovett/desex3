magic
tech c035u
timestamp 1385075154
<< nwell >>
rect 202 526 1443 738
rect 202 524 1332 526
rect 202 493 1331 524
rect 202 492 1318 493
rect 202 490 644 492
rect 352 400 644 490
rect 689 400 981 492
rect 1026 400 1318 492
rect 405 399 451 400
rect 742 399 788 400
rect 1079 399 1125 400
<< polysilicon >>
rect 538 690 545 698
rect 565 690 572 698
rect 592 690 599 698
rect 619 690 626 698
rect 875 690 882 698
rect 902 690 909 698
rect 929 690 936 698
rect 956 690 963 698
rect 1212 690 1219 698
rect 1239 690 1246 698
rect 1266 690 1273 698
rect 1293 690 1300 698
rect 480 612 487 620
rect 507 612 514 620
rect 425 557 432 565
rect 370 458 377 466
rect 817 612 824 620
rect 844 612 851 620
rect 762 557 769 565
rect 707 458 714 466
rect 1154 612 1161 620
rect 1181 612 1188 620
rect 1099 557 1106 565
rect 1044 458 1051 466
rect 1394 639 1396 655
rect 1389 594 1396 639
rect 1389 498 1396 546
rect 1389 460 1396 468
rect 370 386 377 400
rect 425 386 432 400
rect 480 387 487 400
rect 375 370 377 386
rect 430 370 432 386
rect 485 383 487 387
rect 507 383 514 400
rect 538 387 545 400
rect 485 376 514 383
rect 485 371 487 376
rect 543 383 545 387
rect 565 383 572 400
rect 592 383 599 400
rect 619 383 626 400
rect 707 386 714 400
rect 762 386 769 400
rect 817 387 824 400
rect 543 376 626 383
rect 543 371 545 376
rect 370 360 377 370
rect 425 360 432 370
rect 480 360 487 371
rect 538 360 545 371
rect 565 360 572 376
rect 712 370 714 386
rect 767 370 769 386
rect 822 383 824 387
rect 844 383 851 400
rect 875 387 882 400
rect 822 376 851 383
rect 822 371 824 376
rect 880 383 882 387
rect 902 383 909 400
rect 929 383 936 400
rect 956 383 963 400
rect 1044 386 1051 400
rect 1099 386 1106 400
rect 1154 387 1161 400
rect 880 376 963 383
rect 880 371 882 376
rect 707 360 714 370
rect 762 360 769 370
rect 817 360 824 371
rect 875 360 882 371
rect 902 360 909 376
rect 1049 370 1051 386
rect 1104 370 1106 386
rect 1159 383 1161 387
rect 1181 383 1188 400
rect 1212 387 1219 400
rect 1159 376 1188 383
rect 1159 371 1161 376
rect 1217 383 1219 387
rect 1239 383 1246 400
rect 1266 383 1273 400
rect 1293 383 1300 400
rect 1217 376 1300 383
rect 1217 371 1219 376
rect 1044 360 1051 370
rect 1099 360 1106 370
rect 1154 360 1161 371
rect 1212 360 1219 371
rect 1239 360 1246 376
rect 370 332 377 340
rect 425 298 432 306
rect 480 206 487 214
rect 707 332 714 340
rect 762 298 769 306
rect 817 206 824 214
rect 1044 332 1051 340
rect 1099 298 1106 306
rect 1154 206 1161 214
rect 538 152 545 160
rect 565 152 572 160
rect 875 152 882 160
rect 902 152 909 160
rect 1212 152 1219 160
rect 1239 152 1246 160
<< ndiffusion >>
rect 1387 468 1389 498
rect 1396 468 1398 498
rect 368 340 370 360
rect 377 340 379 360
rect 423 306 425 360
rect 432 306 434 360
rect 478 214 480 360
rect 487 214 489 360
rect 536 160 538 360
rect 545 160 547 360
rect 563 160 565 360
rect 572 160 574 360
rect 705 340 707 360
rect 714 340 716 360
rect 760 306 762 360
rect 769 306 771 360
rect 815 214 817 360
rect 824 214 826 360
rect 873 160 875 360
rect 882 160 884 360
rect 900 160 902 360
rect 909 160 911 360
rect 1042 340 1044 360
rect 1051 340 1053 360
rect 1097 306 1099 360
rect 1106 306 1108 360
rect 1152 214 1154 360
rect 1161 214 1163 360
rect 1210 160 1212 360
rect 1219 160 1221 360
rect 1237 160 1239 360
rect 1246 160 1248 360
<< pdiffusion >>
rect 368 400 370 458
rect 377 400 379 458
rect 423 400 425 557
rect 432 400 434 557
rect 478 400 480 612
rect 487 400 489 612
rect 505 400 507 612
rect 514 400 516 612
rect 536 400 538 690
rect 545 400 547 690
rect 563 400 565 690
rect 572 400 574 690
rect 590 400 592 690
rect 599 400 601 690
rect 617 400 619 690
rect 626 400 628 690
rect 705 400 707 458
rect 714 400 716 458
rect 760 400 762 557
rect 769 400 771 557
rect 815 400 817 612
rect 824 400 826 612
rect 842 400 844 612
rect 851 400 853 612
rect 873 400 875 690
rect 882 400 884 690
rect 900 400 902 690
rect 909 400 911 690
rect 927 400 929 690
rect 936 400 938 690
rect 954 400 956 690
rect 963 400 965 690
rect 1042 400 1044 458
rect 1051 400 1053 458
rect 1097 400 1099 557
rect 1106 400 1108 557
rect 1152 400 1154 612
rect 1161 400 1163 612
rect 1179 400 1181 612
rect 1188 400 1190 612
rect 1210 400 1212 690
rect 1219 400 1221 690
rect 1237 400 1239 690
rect 1246 400 1248 690
rect 1264 400 1266 690
rect 1273 400 1275 690
rect 1291 400 1293 690
rect 1300 400 1302 690
rect 1387 546 1389 594
rect 1396 546 1398 594
<< pohmic >>
rect 320 78 326 88
rect 342 78 354 88
rect 370 78 382 88
rect 398 78 410 88
rect 426 78 438 88
rect 454 78 466 88
rect 482 78 494 88
rect 510 78 522 88
rect 538 78 550 88
rect 567 78 579 88
rect 595 78 607 88
rect 623 78 635 88
rect 651 78 663 88
rect 679 78 691 88
rect 707 78 719 88
rect 735 78 747 88
rect 763 78 775 88
rect 791 78 803 88
rect 819 78 831 88
rect 847 78 859 88
rect 875 78 887 88
rect 904 78 916 88
rect 932 78 944 88
rect 960 78 972 88
rect 988 78 1000 88
rect 1016 78 1028 88
rect 1044 78 1056 88
rect 1072 78 1084 88
rect 1100 78 1112 88
rect 1128 78 1140 88
rect 1156 78 1168 88
rect 1184 78 1196 88
rect 1212 78 1224 88
rect 1241 78 1253 88
rect 1269 78 1281 88
rect 1297 78 1309 88
rect 1325 78 1337 88
rect 1353 78 1365 88
rect 1381 78 1393 88
rect 1409 78 1421 88
rect 1437 78 1443 88
<< nohmic >>
rect 202 728 214 738
rect 230 728 242 738
rect 258 728 270 738
rect 286 728 298 738
rect 314 728 326 738
rect 342 728 354 738
rect 370 728 382 738
rect 398 728 410 738
rect 426 728 438 738
rect 454 728 466 738
rect 482 728 494 738
rect 510 728 522 738
rect 538 728 550 738
rect 567 728 579 738
rect 595 728 607 738
rect 623 728 635 738
rect 651 728 663 738
rect 679 728 691 738
rect 707 728 719 738
rect 735 728 747 738
rect 763 728 775 738
rect 791 728 803 738
rect 819 728 831 738
rect 847 728 859 738
rect 875 728 887 738
rect 904 728 916 738
rect 932 728 944 738
rect 960 728 972 738
rect 988 728 1000 738
rect 1016 728 1028 738
rect 1044 728 1056 738
rect 1072 728 1084 738
rect 1100 728 1112 738
rect 1128 728 1140 738
rect 1156 728 1168 738
rect 1184 728 1196 738
rect 1212 728 1224 738
rect 1241 728 1253 738
rect 1269 728 1281 738
rect 1297 728 1309 738
rect 1325 728 1337 738
rect 1353 728 1365 738
rect 1381 728 1393 738
rect 1409 728 1421 738
rect 1437 728 1443 738
<< ntransistor >>
rect 1389 468 1396 498
rect 370 340 377 360
rect 425 306 432 360
rect 480 214 487 360
rect 538 160 545 360
rect 565 160 572 360
rect 707 340 714 360
rect 762 306 769 360
rect 817 214 824 360
rect 875 160 882 360
rect 902 160 909 360
rect 1044 340 1051 360
rect 1099 306 1106 360
rect 1154 214 1161 360
rect 1212 160 1219 360
rect 1239 160 1246 360
<< ptransistor >>
rect 370 400 377 458
rect 425 400 432 557
rect 480 400 487 612
rect 507 400 514 612
rect 538 400 545 690
rect 565 400 572 690
rect 592 400 599 690
rect 619 400 626 690
rect 707 400 714 458
rect 762 400 769 557
rect 817 400 824 612
rect 844 400 851 612
rect 875 400 882 690
rect 902 400 909 690
rect 929 400 936 690
rect 956 400 963 690
rect 1044 400 1051 458
rect 1099 400 1106 557
rect 1154 400 1161 612
rect 1181 400 1188 612
rect 1212 400 1219 690
rect 1239 400 1246 690
rect 1266 400 1273 690
rect 1293 400 1300 690
rect 1389 546 1396 594
<< polycontact >>
rect 1378 639 1394 655
rect 359 370 375 386
rect 414 370 430 386
rect 469 371 485 387
rect 527 371 543 387
rect 696 370 712 386
rect 751 370 767 386
rect 806 371 822 387
rect 864 371 880 387
rect 1033 370 1049 386
rect 1088 370 1104 386
rect 1143 371 1159 387
rect 1201 371 1217 387
<< ndiffcontact >>
rect 1371 468 1387 498
rect 1398 468 1414 498
rect 352 340 368 360
rect 379 340 395 360
rect 407 306 423 360
rect 434 306 450 360
rect 462 214 478 360
rect 489 214 505 360
rect 520 160 536 360
rect 547 160 563 360
rect 574 160 590 360
rect 689 340 705 360
rect 716 340 732 360
rect 744 306 760 360
rect 771 306 787 360
rect 799 214 815 360
rect 826 214 842 360
rect 857 160 873 360
rect 884 160 900 360
rect 911 160 927 360
rect 1026 340 1042 360
rect 1053 340 1069 360
rect 1081 306 1097 360
rect 1108 306 1124 360
rect 1136 214 1152 360
rect 1163 214 1179 360
rect 1194 160 1210 360
rect 1221 160 1237 360
rect 1248 160 1264 360
<< pdiffcontact >>
rect 519 612 536 690
rect 352 400 368 458
rect 379 400 395 458
rect 407 400 423 557
rect 434 400 450 557
rect 462 400 478 612
rect 489 400 505 612
rect 516 400 536 612
rect 547 400 563 690
rect 574 400 590 690
rect 601 400 617 690
rect 628 400 644 690
rect 856 612 873 690
rect 689 400 705 458
rect 716 400 732 458
rect 744 400 760 557
rect 771 400 787 557
rect 799 400 815 612
rect 826 400 842 612
rect 853 400 873 612
rect 884 400 900 690
rect 911 400 927 690
rect 938 400 954 690
rect 965 400 981 690
rect 1193 612 1210 690
rect 1026 400 1042 458
rect 1053 400 1069 458
rect 1081 400 1097 557
rect 1108 400 1124 557
rect 1136 400 1152 612
rect 1163 400 1179 612
rect 1190 400 1210 612
rect 1221 400 1237 690
rect 1248 400 1264 690
rect 1275 400 1291 690
rect 1302 400 1318 690
rect 1371 546 1387 594
rect 1398 546 1414 594
<< psubstratetap >>
rect 326 78 342 94
rect 354 78 370 94
rect 382 78 398 94
rect 410 78 426 94
rect 438 78 454 94
rect 466 78 482 94
rect 494 78 510 94
rect 522 78 538 94
rect 550 78 567 94
rect 579 78 595 94
rect 607 78 623 94
rect 635 78 651 94
rect 663 78 679 94
rect 691 78 707 94
rect 719 78 735 94
rect 747 78 763 94
rect 775 78 791 94
rect 803 78 819 94
rect 831 78 847 94
rect 859 78 875 94
rect 887 78 904 94
rect 916 78 932 94
rect 944 78 960 94
rect 972 78 988 94
rect 1000 78 1016 94
rect 1028 78 1044 94
rect 1056 78 1072 94
rect 1084 78 1100 94
rect 1112 78 1128 94
rect 1140 78 1156 94
rect 1168 78 1184 94
rect 1196 78 1212 94
rect 1224 78 1241 94
rect 1253 78 1269 94
rect 1281 78 1297 94
rect 1309 78 1325 94
rect 1337 78 1353 94
rect 1365 78 1381 94
rect 1393 78 1409 94
rect 1421 78 1437 94
<< nsubstratetap >>
rect 214 722 230 738
rect 242 722 258 738
rect 270 722 286 738
rect 298 722 314 738
rect 326 722 342 738
rect 354 722 370 738
rect 382 722 398 738
rect 410 722 426 738
rect 438 722 454 738
rect 466 722 482 738
rect 494 722 510 738
rect 522 722 538 738
rect 550 722 567 738
rect 579 722 595 738
rect 607 722 623 738
rect 635 722 651 738
rect 663 722 679 738
rect 691 722 707 738
rect 719 722 735 738
rect 747 722 763 738
rect 775 722 791 738
rect 803 722 819 738
rect 831 722 847 738
rect 859 722 875 738
rect 887 722 904 738
rect 916 722 932 738
rect 944 722 960 738
rect 972 722 988 738
rect 1000 722 1016 738
rect 1028 722 1044 738
rect 1056 722 1072 738
rect 1084 722 1100 738
rect 1112 722 1128 738
rect 1140 722 1156 738
rect 1168 722 1184 738
rect 1196 722 1212 738
rect 1224 722 1241 738
rect 1253 722 1269 738
rect 1281 722 1297 738
rect 1309 722 1325 738
rect 1337 722 1353 738
rect 1365 722 1381 738
rect 1393 722 1409 738
rect 1421 722 1437 738
<< metal1 >>
rect 236 774 1356 784
rect 1400 774 1443 784
rect 236 751 1443 761
rect 200 722 214 738
rect 230 722 242 738
rect 258 722 270 738
rect 286 722 298 738
rect 314 722 326 738
rect 342 722 354 738
rect 370 722 382 738
rect 398 722 410 738
rect 426 722 438 738
rect 454 722 466 738
rect 482 722 494 738
rect 510 722 522 738
rect 538 722 550 738
rect 567 722 579 738
rect 595 722 607 738
rect 623 722 635 738
rect 651 722 663 738
rect 679 722 691 738
rect 707 722 719 738
rect 735 722 747 738
rect 763 722 775 738
rect 791 722 803 738
rect 819 722 831 738
rect 847 722 859 738
rect 875 722 887 738
rect 904 722 916 738
rect 932 722 944 738
rect 960 722 972 738
rect 988 722 1000 738
rect 1016 722 1028 738
rect 1044 722 1056 738
rect 1072 722 1084 738
rect 1100 722 1112 738
rect 1128 722 1140 738
rect 1156 722 1168 738
rect 1184 722 1196 738
rect 1212 722 1224 738
rect 1241 722 1253 738
rect 1269 722 1281 738
rect 1297 722 1309 738
rect 1325 722 1337 738
rect 1353 722 1365 738
rect 1381 722 1393 738
rect 1409 722 1421 738
rect 1437 722 1443 738
rect 200 713 1443 722
rect 352 458 368 713
rect 407 557 423 713
rect 462 612 478 713
rect 516 690 536 713
rect 574 690 590 713
rect 628 690 644 713
rect 516 612 519 690
rect 689 458 705 713
rect 744 557 760 713
rect 799 612 815 713
rect 853 690 873 713
rect 911 690 927 713
rect 965 690 981 713
rect 853 612 856 690
rect 1026 458 1042 713
rect 1081 557 1097 713
rect 1136 612 1152 713
rect 1190 690 1210 713
rect 1248 690 1264 713
rect 1302 690 1318 713
rect 1190 612 1193 690
rect 1380 655 1394 661
rect 1404 594 1414 713
rect 1371 498 1381 546
rect 284 373 359 383
rect 385 383 395 400
rect 385 373 414 383
rect 385 360 395 373
rect 440 384 450 400
rect 440 374 469 384
rect 440 360 450 374
rect 495 384 505 400
rect 495 374 527 384
rect 495 360 505 374
rect 553 385 563 400
rect 607 387 617 400
rect 553 375 606 385
rect 553 360 563 375
rect 667 373 696 383
rect 722 383 732 400
rect 722 373 751 383
rect 722 360 732 373
rect 777 384 787 400
rect 777 374 806 384
rect 777 360 787 374
rect 832 384 842 400
rect 832 374 864 384
rect 832 360 842 374
rect 890 385 900 400
rect 944 387 954 400
rect 890 375 944 385
rect 890 360 900 375
rect 1022 373 1033 383
rect 1059 383 1069 400
rect 1059 373 1088 383
rect 1059 360 1069 373
rect 1114 384 1124 400
rect 1114 374 1143 384
rect 1114 360 1124 374
rect 1169 384 1179 400
rect 1169 374 1201 384
rect 1169 360 1179 374
rect 1227 385 1237 400
rect 1281 387 1291 400
rect 1227 375 1279 385
rect 1227 360 1237 375
rect 352 103 368 340
rect 407 103 423 306
rect 462 103 478 214
rect 520 103 536 160
rect 574 103 590 160
rect 689 103 705 340
rect 744 103 760 306
rect 799 103 815 214
rect 857 103 873 160
rect 911 103 927 160
rect 1026 103 1042 340
rect 1081 103 1097 306
rect 1136 103 1152 214
rect 1194 103 1210 160
rect 1248 103 1264 160
rect 1398 103 1408 468
rect 320 94 1443 103
rect 320 78 326 94
rect 342 78 354 94
rect 370 78 382 94
rect 398 78 410 94
rect 426 78 438 94
rect 454 78 466 94
rect 482 78 494 94
rect 510 78 522 94
rect 538 78 550 94
rect 567 78 579 94
rect 595 78 607 94
rect 623 78 635 94
rect 651 78 663 94
rect 679 78 691 94
rect 707 78 719 94
rect 735 78 747 94
rect 763 78 775 94
rect 791 78 803 94
rect 819 78 831 94
rect 847 78 859 94
rect 875 78 887 94
rect 904 78 916 94
rect 932 78 944 94
rect 960 78 972 94
rect 988 78 1000 94
rect 1016 78 1028 94
rect 1044 78 1056 94
rect 1072 78 1084 94
rect 1100 78 1112 94
rect 1128 78 1140 94
rect 1156 78 1168 94
rect 1184 78 1196 94
rect 1212 78 1224 94
rect 1241 78 1253 94
rect 1269 78 1281 94
rect 1297 78 1309 94
rect 1325 78 1337 94
rect 1353 78 1365 94
rect 1381 78 1393 94
rect 1409 78 1421 94
rect 1437 78 1443 94
rect 620 55 1443 65
rect 260 32 653 42
rect 959 32 1443 42
rect 308 9 1009 19
rect 1294 9 1443 19
<< m2contact >>
rect 222 773 236 787
rect 1356 773 1370 787
rect 1386 773 1400 787
rect 222 749 236 763
rect 0 713 200 738
rect 1380 661 1394 675
rect 1357 580 1371 594
rect 270 371 284 385
rect 606 373 620 387
rect 653 371 667 385
rect 944 373 958 387
rect 1008 371 1022 385
rect 1279 373 1293 387
rect 606 53 620 67
rect 246 29 260 43
rect 653 30 667 44
rect 945 31 959 45
rect 294 5 308 19
rect 1009 7 1023 21
rect 1280 7 1294 21
<< metal2 >>
rect 0 738 200 792
rect 223 787 235 792
rect 0 0 200 713
rect 223 0 235 749
rect 247 43 259 792
rect 271 385 283 792
rect 247 0 259 29
rect 271 0 283 371
rect 295 19 307 792
rect 1358 594 1370 773
rect 1386 675 1398 773
rect 1394 661 1398 675
rect 607 67 619 373
rect 654 44 666 371
rect 946 45 958 373
rect 1010 21 1022 371
rect 1281 21 1293 373
rect 295 0 307 5
<< labels >>
rlabel metal2 0 792 200 792 5 Vdd!
rlabel metal2 223 792 235 792 5 SDO
rlabel metal2 247 792 259 792 5 Test
rlabel metal2 271 792 283 792 5 Clock
rlabel metal2 295 792 307 792 5 nReset
rlabel metal2 247 0 259 0 1 Test
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 295 0 307 0 1 nReset
rlabel metal2 223 0 235 0 1 SDI
rlabel metal1 1443 713 1443 738 7 Vdd!
rlabel metal1 1443 751 1443 761 7 SDI
rlabel metal1 1443 774 1443 784 7 nSDO
rlabel metal1 1443 55 1443 65 7 ClockOut
rlabel metal1 1443 32 1443 42 7 TestOut
rlabel metal1 1443 9 1443 19 7 nResetOut
rlabel metal1 1443 78 1443 103 7 GND!
<< end >>
