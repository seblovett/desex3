magic
tech c035u
timestamp 1385631125
<< nwell >>
rect 0 408 264 752
<< polysilicon >>
rect 24 691 31 699
rect 51 691 58 717
rect 147 691 154 699
rect 177 691 184 699
rect 232 691 239 699
rect 24 613 31 643
rect 51 613 58 643
rect 106 613 113 659
rect 24 192 31 565
rect 51 192 58 565
rect 106 192 113 565
rect 147 555 154 643
rect 177 613 184 643
rect 232 583 239 643
rect 238 567 239 583
rect 147 218 154 539
rect 177 270 184 565
rect 24 132 31 162
rect 51 132 58 162
rect 106 152 113 162
rect 147 132 154 202
rect 177 192 184 254
rect 232 208 239 567
rect 177 132 184 162
rect 232 132 239 192
rect 24 94 31 102
rect 51 94 58 102
rect 147 94 154 102
rect 177 94 184 102
rect 232 94 239 102
<< ndiffusion >>
rect 22 162 24 192
rect 31 162 51 192
rect 58 162 60 192
rect 104 162 106 192
rect 113 162 115 192
rect 175 162 177 192
rect 184 162 186 192
rect 22 102 24 132
rect 31 102 33 132
rect 49 102 51 132
rect 58 102 60 132
rect 145 102 147 132
rect 154 102 177 132
rect 184 102 186 132
rect 230 102 232 132
rect 239 102 241 132
<< pdiffusion >>
rect 22 643 24 691
rect 31 643 51 691
rect 58 643 60 691
rect 145 643 147 691
rect 154 643 159 691
rect 175 643 177 691
rect 184 643 186 691
rect 202 643 232 691
rect 239 643 241 691
rect 22 565 24 613
rect 31 565 33 613
rect 49 565 51 613
rect 58 565 60 613
rect 76 565 106 613
rect 113 565 115 613
rect 175 565 177 613
rect 184 565 186 613
<< pohmic >>
rect 0 67 6 77
rect 22 67 34 77
rect 50 67 62 77
rect 78 67 90 77
rect 106 67 118 77
rect 134 67 146 77
rect 162 67 174 77
rect 190 67 202 77
rect 218 67 230 77
rect 246 67 264 77
<< nohmic >>
rect 0 742 6 752
rect 22 742 34 752
rect 50 742 62 752
rect 78 742 90 752
rect 106 742 118 752
rect 134 742 146 752
rect 162 742 174 752
rect 190 742 202 752
rect 218 742 230 752
rect 246 742 264 752
<< ntransistor >>
rect 24 162 31 192
rect 51 162 58 192
rect 106 162 113 192
rect 177 162 184 192
rect 24 102 31 132
rect 51 102 58 132
rect 147 102 154 132
rect 177 102 184 132
rect 232 102 239 132
<< ptransistor >>
rect 24 643 31 691
rect 51 643 58 691
rect 147 643 154 691
rect 177 643 184 691
rect 232 643 239 691
rect 24 565 31 613
rect 51 565 58 613
rect 106 565 113 613
rect 177 565 184 613
<< polycontact >>
rect 101 659 117 675
rect 222 567 238 583
rect 138 539 154 555
rect 168 254 184 270
rect 138 202 154 218
rect 101 136 117 152
rect 223 192 239 208
<< ndiffcontact >>
rect 6 162 22 192
rect 60 162 76 192
rect 88 162 104 192
rect 115 162 131 192
rect 159 162 175 192
rect 186 162 202 192
rect 6 102 22 132
rect 33 102 49 132
rect 60 102 76 132
rect 129 102 145 132
rect 186 102 202 132
rect 214 102 230 132
rect 241 102 257 132
<< pdiffcontact >>
rect 6 643 22 691
rect 60 643 76 691
rect 129 643 145 691
rect 159 643 175 691
rect 186 643 202 691
rect 241 643 257 691
rect 6 565 22 613
rect 33 565 49 613
rect 60 565 76 613
rect 115 565 131 613
rect 159 565 175 613
rect 186 565 202 613
<< psubstratetap >>
rect 6 67 22 83
rect 34 67 50 83
rect 62 67 78 83
rect 90 67 106 83
rect 118 67 134 83
rect 146 67 162 83
rect 174 67 190 83
rect 202 67 218 83
rect 230 67 246 83
<< nsubstratetap >>
rect 6 736 22 752
rect 34 736 50 752
rect 62 736 78 752
rect 90 736 106 752
rect 118 736 134 752
rect 146 736 162 752
rect 174 736 190 752
rect 202 736 218 752
rect 230 736 246 752
<< metal1 >>
rect 0 782 264 792
rect 0 762 264 772
rect 0 736 6 752
rect 22 736 34 752
rect 50 736 62 752
rect 78 736 90 752
rect 106 736 118 752
rect 134 736 146 752
rect 162 736 174 752
rect 190 736 202 752
rect 218 736 230 752
rect 246 736 264 752
rect 0 727 264 736
rect 9 691 19 727
rect 132 691 142 727
rect 189 691 199 727
rect 76 662 101 672
rect 9 633 19 643
rect 135 633 145 643
rect 162 633 172 643
rect 9 623 73 633
rect 135 623 152 633
rect 162 623 231 633
rect 9 613 19 623
rect 63 613 73 623
rect 142 613 152 623
rect 142 603 159 613
rect 221 583 231 623
rect 243 607 253 643
rect 221 567 222 583
rect 36 267 46 565
rect 118 552 128 565
rect 192 555 202 565
rect 118 541 138 552
rect 36 257 168 267
rect 63 192 73 257
rect 91 208 138 218
rect 91 192 101 208
rect 192 192 202 218
rect 131 172 159 182
rect 9 132 19 162
rect 36 142 101 152
rect 36 132 46 142
rect 131 132 141 172
rect 222 192 223 208
rect 222 152 232 192
rect 189 142 232 152
rect 189 132 199 142
rect 244 132 254 168
rect 9 92 19 102
rect 63 92 73 102
rect 132 92 142 102
rect 217 92 227 102
rect 0 83 264 92
rect 0 67 6 83
rect 22 67 34 83
rect 50 67 62 83
rect 78 67 90 83
rect 106 67 118 83
rect 134 67 146 83
rect 162 67 174 83
rect 190 67 202 83
rect 218 67 230 83
rect 246 67 264 83
rect 0 47 264 57
rect 0 27 264 37
rect 0 7 264 17
<< m2contact >>
rect 47 703 61 717
rect 241 593 255 607
rect 191 541 205 555
rect 24 208 38 222
rect 191 218 205 232
rect 242 168 256 182
<< metal2 >>
rect 24 222 36 799
rect 48 717 60 799
rect 24 0 36 208
rect 48 0 60 703
rect 192 555 204 799
rect 240 607 252 799
rect 240 593 241 607
rect 192 232 204 541
rect 192 0 204 218
rect 240 182 252 593
rect 240 168 242 182
rect 240 0 252 168
<< labels >>
rlabel metal1 0 67 0 92 3 GND!
rlabel metal1 0 47 0 57 3 Clock
rlabel metal1 0 27 0 37 3 Test
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 727 0 752 3 Vdd!
rlabel metal1 264 27 264 37 7 Test
rlabel metal1 264 47 264 57 7 Clock
rlabel metal1 264 67 264 92 7 GND!
rlabel metal1 264 727 264 752 7 Vdd!
rlabel metal1 264 782 264 792 7 ScanReturn
rlabel metal2 240 799 252 799 5 S
rlabel metal2 192 799 204 799 5 C
rlabel metal2 48 799 60 799 5 B
rlabel metal2 24 799 36 799 5 A
rlabel metal2 24 0 36 0 1 A
rlabel metal2 48 0 60 0 1 B
rlabel metal2 192 0 204 0 1 C
rlabel metal2 240 0 252 0 1 S
rlabel metal1 0 762 0 772 3 Scan
rlabel metal1 264 762 264 772 7 Scan
rlabel metal1 0 7 0 17 3 nReset
rlabel metal1 264 7 264 17 7 nReset
<< end >>
