magic
tech c035u
timestamp 1386235218
<< nwell >>
rect 0 401 192 799
<< pwell >>
rect 0 0 192 401
<< polysilicon >>
rect 34 691 41 699
rect 64 691 71 699
rect 91 691 98 699
rect 118 691 125 699
rect 149 691 156 699
rect 34 612 41 643
rect 64 599 71 643
rect 34 485 41 564
rect 34 347 41 469
rect 64 347 71 583
rect 91 500 98 643
rect 118 488 125 643
rect 149 633 156 643
rect 152 617 156 633
rect 91 347 98 484
rect 118 347 125 472
rect 149 393 156 617
rect 151 377 156 393
rect 34 282 41 317
rect 64 278 71 317
rect 91 309 98 317
rect 118 309 125 317
rect 149 282 156 377
rect 34 243 41 252
rect 149 244 156 252
<< ndiffusion >>
rect 32 317 34 347
rect 41 317 43 347
rect 59 317 64 347
rect 71 317 91 347
rect 98 317 100 347
rect 116 317 118 347
rect 125 317 127 347
rect 32 252 34 282
rect 41 252 43 282
rect 147 252 149 282
rect 156 252 158 282
<< pdiffusion >>
rect 32 643 34 691
rect 41 643 43 691
rect 59 643 64 691
rect 71 643 73 691
rect 89 643 91 691
rect 98 643 100 691
rect 116 643 118 691
rect 125 643 128 691
rect 144 643 149 691
rect 156 643 159 691
rect 32 564 34 612
rect 41 564 43 612
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 192 86
rect 0 76 192 79
<< nohmic >>
rect 0 743 192 746
rect 0 736 8 743
rect 24 736 36 743
rect 52 736 64 743
rect 80 736 92 743
rect 108 736 121 743
rect 137 736 149 743
rect 165 736 192 743
<< ntransistor >>
rect 34 317 41 347
rect 64 317 71 347
rect 91 317 98 347
rect 118 317 125 347
rect 34 252 41 282
rect 149 252 156 282
<< ptransistor >>
rect 34 643 41 691
rect 64 643 71 691
rect 91 643 98 691
rect 118 643 125 691
rect 149 643 156 691
rect 34 564 41 612
<< polycontact >>
rect 64 583 80 599
rect 30 469 46 485
rect 84 484 100 500
rect 136 617 152 633
rect 118 472 134 488
rect 135 377 151 393
rect 64 262 80 278
<< ndiffcontact >>
rect 16 317 32 347
rect 43 317 59 347
rect 100 317 116 347
rect 127 317 143 347
rect 16 252 32 282
rect 43 252 59 282
rect 131 252 147 282
rect 158 252 174 282
<< pdiffcontact >>
rect 16 643 32 691
rect 43 643 59 691
rect 73 643 89 691
rect 100 643 116 691
rect 128 643 144 691
rect 159 643 175 691
rect 16 564 32 612
rect 43 564 59 612
<< psubstratetap >>
rect 100 238 116 254
rect 6 79 22 95
rect 34 79 50 95
rect 62 79 78 95
rect 90 79 106 95
rect 118 79 134 95
rect 146 79 162 95
<< nsubstratetap >>
rect 8 727 24 743
rect 36 727 52 743
rect 64 727 80 743
rect 92 727 108 743
rect 121 727 137 743
rect 149 727 165 743
<< metal1 >>
rect 0 782 192 792
rect 0 759 192 769
rect 0 743 192 746
rect 0 727 8 743
rect 24 727 36 743
rect 52 727 64 743
rect 80 727 92 743
rect 108 727 121 743
rect 137 727 149 743
rect 165 727 192 743
rect 0 721 192 727
rect 16 691 32 721
rect 46 701 113 711
rect 46 691 56 701
rect 103 691 113 701
rect 128 691 144 721
rect 16 612 32 643
rect 76 629 86 643
rect 76 619 136 629
rect 59 583 64 599
rect 162 469 172 643
rect 165 455 172 469
rect 46 380 135 390
rect 46 347 56 380
rect 78 357 140 367
rect 19 307 29 317
rect 78 307 88 357
rect 130 347 140 357
rect 19 297 88 307
rect 100 282 116 317
rect 162 282 172 455
rect 59 262 64 278
rect 100 254 131 282
rect 16 101 32 252
rect 116 252 131 254
rect 100 101 116 238
rect 0 95 192 101
rect 0 79 6 95
rect 22 79 34 95
rect 50 79 62 95
rect 78 79 90 95
rect 106 79 118 95
rect 134 79 146 95
rect 162 79 192 95
rect 0 76 192 79
rect 0 53 192 63
rect 0 30 192 40
rect 0 7 192 17
<< m2contact >>
rect 70 485 84 499
rect 119 488 133 502
rect 46 470 60 484
rect 151 455 165 469
<< metal2 >>
rect 48 484 60 799
rect 72 499 84 799
rect 120 502 132 799
rect 48 0 60 470
rect 72 0 84 485
rect 120 0 132 488
rect 144 469 156 799
rect 144 455 151 469
rect 144 0 156 455
<< labels >>
rlabel metal1 0 76 0 101 1 GND!
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 3 Clock
rlabel metal2 48 0 60 0 1 S
rlabel metal2 144 0 156 0 1 Y
rlabel metal2 72 0 84 0 1 I0
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal2 48 799 60 799 5 S
rlabel metal2 144 799 156 799 5 Y
rlabel metal2 120 799 132 799 5 I1
rlabel metal2 72 799 84 799 5 I0
rlabel metal1 192 76 192 101 7 GND!
rlabel metal1 192 7 192 17 8 nReset
rlabel metal1 192 30 192 40 7 Test
rlabel metal1 192 53 192 63 7 Clock
rlabel metal1 192 721 192 746 7 Vdd!
rlabel metal1 192 782 192 792 6 ScanReturn
rlabel metal1 192 759 192 769 7 Scan
rlabel metal2 120 0 132 0 1 I1
<< end >>
