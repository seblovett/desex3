magic
tech c035u
timestamp 1385634731
<< metal1 >>
rect 236 908 2680 918
rect 2694 908 2800 918
rect 2814 908 2920 918
rect 1464 865 1577 875
rect 3017 865 3097 875
rect 1464 842 1577 852
rect 3017 842 3097 852
rect 1464 804 1577 829
rect 3017 804 3097 829
rect 1464 159 1577 184
rect 3017 159 3097 184
rect 1464 136 1529 146
rect 1543 136 1577 146
rect 3017 136 3097 146
rect 1464 113 1506 123
rect 1520 113 1577 123
rect 3017 113 3097 123
rect 1464 90 1482 100
rect 1496 90 1577 100
rect 3017 90 3097 100
rect 1543 50 1600 60
rect 1614 50 1720 60
rect 1734 50 1840 60
rect 1520 28 1960 38
rect 1974 28 2080 38
rect 2094 28 2200 38
rect 1497 4 2320 14
rect 2334 4 2440 14
rect 2454 4 2560 14
<< m2contact >>
rect 222 907 236 921
rect 2680 906 2694 920
rect 2800 906 2814 920
rect 2920 906 2934 920
rect 1529 134 1543 148
rect 1506 110 1520 124
rect 1482 87 1496 101
rect 1529 50 1543 64
rect 1600 48 1614 62
rect 1720 48 1734 62
rect 1840 48 1854 62
rect 1506 26 1520 40
rect 1960 26 1974 40
rect 2080 26 2094 40
rect 2200 26 2214 40
rect 1483 2 1497 16
rect 2320 2 2334 16
rect 2440 2 2454 16
rect 2560 2 2574 16
<< metal2 >>
rect 223 921 235 934
rect 223 882 235 907
rect 2681 882 2693 906
rect 2801 882 2813 906
rect 2921 882 2933 906
rect 0 0 200 83
rect 223 0 235 83
rect 247 0 259 83
rect 271 0 283 83
rect 295 0 307 83
rect 1484 16 1496 87
rect 1507 40 1519 110
rect 1530 64 1542 134
rect 1601 62 1613 83
rect 1721 62 1733 83
rect 1841 62 1853 83
rect 1961 40 1973 83
rect 2081 40 2093 83
rect 2201 40 2213 83
rect 2321 16 2333 83
rect 2441 16 2453 83
rect 2561 16 2573 83
use leftbuf leftbuf_0
timestamp 1385634621
transform 1 0 0 0 1 93
box 0 -10 1464 789
use inv inv_0
timestamp 1385631115
transform 1 0 1577 0 1 83
box 0 0 120 799
use inv inv_1
timestamp 1385631115
transform 1 0 1697 0 1 83
box 0 0 120 799
use inv inv_2
timestamp 1385631115
transform 1 0 1817 0 1 83
box 0 0 120 799
use inv inv_3
timestamp 1385631115
transform 1 0 1937 0 1 83
box 0 0 120 799
use inv inv_4
timestamp 1385631115
transform 1 0 2057 0 1 83
box 0 0 120 799
use inv inv_5
timestamp 1385631115
transform 1 0 2177 0 1 83
box 0 0 120 799
use inv inv_6
timestamp 1385631115
transform 1 0 2297 0 1 83
box 0 0 120 799
use inv inv_7
timestamp 1385631115
transform 1 0 2417 0 1 83
box 0 0 120 799
use inv inv_8
timestamp 1385631115
transform 1 0 2537 0 1 83
box 0 0 120 799
use inv inv_9
timestamp 1385631115
transform 1 0 2657 0 1 83
box 0 0 120 799
use inv inv_10
timestamp 1385631115
transform 1 0 2777 0 1 83
box 0 0 120 799
use inv inv_11
timestamp 1385631115
transform 1 0 2897 0 1 83
box 0 0 120 799
<< labels >>
rlabel metal2 223 934 235 934 5 SDO
rlabel metal2 295 0 307 0 1 nReset
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 247 0 259 0 1 Test
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal1 3097 159 3097 184 7 GND!
rlabel metal1 3097 136 3097 146 7 ClockOut
rlabel metal1 3097 113 3097 123 7 TestOut
rlabel metal1 3097 90 3097 100 7 nResetOut
rlabel metal1 3097 804 3097 829 7 Vdd!
rlabel metal1 3097 842 3097 852 7 SDI
rlabel metal1 3097 865 3097 875 7 nSDO
<< end >>
