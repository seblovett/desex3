magic
tech c035u
timestamp 1385998521
<< nwell >>
rect 0 402 96 746
<< polysilicon >>
rect 28 595 35 603
rect 55 595 62 603
rect 28 365 35 547
rect 55 427 62 547
rect 61 411 62 427
rect 28 339 35 349
rect 55 339 62 411
rect 28 301 35 309
rect 55 301 62 309
<< ndiffusion >>
rect 26 309 28 339
rect 35 309 55 339
rect 62 309 64 339
<< pdiffusion >>
rect 26 547 28 595
rect 35 547 37 595
rect 53 547 55 595
rect 62 547 64 595
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 96 86
rect 0 76 96 79
<< nohmic >>
rect 0 743 96 746
rect 0 736 6 743
rect 22 736 34 743
rect 50 736 62 743
rect 78 736 96 743
<< ntransistor >>
rect 28 309 35 339
rect 55 309 62 339
<< ptransistor >>
rect 28 547 35 595
rect 55 547 62 595
<< polycontact >>
rect 45 411 61 427
rect 24 349 40 365
<< ndiffcontact >>
rect 10 309 26 339
rect 64 309 80 339
<< pdiffcontact >>
rect 10 547 26 595
rect 37 547 53 595
rect 64 547 80 595
<< psubstratetap >>
rect 6 79 22 95
rect 34 79 50 95
rect 62 79 78 95
<< nsubstratetap >>
rect 6 727 22 743
rect 34 727 50 743
rect 62 727 78 743
<< metal1 >>
rect 0 782 96 792
rect 0 759 96 769
rect 0 743 96 746
rect 0 727 6 743
rect 22 727 34 743
rect 50 727 62 743
rect 78 727 96 743
rect 0 721 96 727
rect 10 595 26 721
rect 64 595 80 721
rect 37 487 47 547
rect 37 477 71 487
rect 71 401 81 473
rect 70 391 81 401
rect 70 339 80 391
rect 10 101 26 309
rect 0 95 96 101
rect 0 79 6 95
rect 22 79 34 95
rect 50 79 62 95
rect 78 79 96 95
rect 0 76 96 79
rect 0 53 96 63
rect 0 30 96 40
rect 0 7 96 17
<< m2contact >>
rect 71 473 85 487
rect 46 397 60 411
rect 24 365 38 379
<< metal2 >>
rect 24 722 36 799
rect 23 595 36 722
rect 24 547 37 595
rect 24 379 36 547
rect 48 427 60 799
rect 72 487 84 799
rect 48 411 61 427
rect 24 349 38 365
rect 24 0 36 349
rect 48 0 60 397
rect 72 95 84 473
rect 71 79 84 95
rect 72 0 84 79
<< labels >>
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 96 53 96 63 7 Clock
rlabel metal1 96 30 96 40 7 Test
rlabel metal1 96 7 96 17 8 nReset
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 96 721 96 746 7 Vdd!
rlabel metal1 96 759 96 769 7 Scan
rlabel metal1 96 782 96 792 6 ScanReturn
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal2 72 0 84 0 1 Y
rlabel metal2 48 0 60 0 1 B
rlabel metal2 24 0 36 0 1 A
rlabel metal2 72 799 84 799 5 Y
rlabel metal2 48 799 60 799 5 B
rlabel metal2 24 799 36 799 5 A
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 96 76 96 101 7 GND!
<< end >>
