magic
tech c035u
timestamp 1384718636
<< error_p >>
rect 222 90 229 97
<< nwell >>
rect 18 310 358 610
rect 19 298 358 310
rect 19 240 359 298
<< polysilicon >>
rect 37 436 44 506
rect 71 496 78 543
rect 106 496 113 579
rect 186 501 229 508
rect 186 496 193 501
rect 222 496 229 501
rect 260 496 267 610
rect 333 496 340 610
rect 37 80 44 388
rect 71 352 78 448
rect 106 436 113 448
rect 145 436 152 444
rect 186 436 193 446
rect 222 436 229 448
rect 106 352 113 388
rect 145 352 152 388
rect 186 352 193 388
rect 222 352 229 388
rect 260 378 267 448
rect 333 436 340 480
rect 71 146 78 304
rect 106 198 113 304
rect 145 294 152 304
rect 145 198 152 278
rect 106 146 113 168
rect 37 1 44 50
rect 71 38 78 116
rect 106 80 113 116
rect 145 80 152 168
rect 186 146 193 304
rect 222 294 229 304
rect 222 146 229 278
rect 186 66 193 116
rect 222 106 229 116
rect 222 80 229 90
rect 260 80 267 362
rect 292 352 299 388
rect 292 172 299 304
rect 333 198 340 388
rect 292 146 299 156
rect 71 0 78 8
rect 106 1 113 50
rect 145 18 152 50
rect 186 38 193 50
rect 222 38 229 50
rect 260 39 267 50
rect 186 0 193 8
rect 222 0 229 8
rect 260 1 267 8
rect 292 1 299 116
rect 333 80 340 168
rect 333 1 340 50
<< ndiffusion >>
rect 104 168 106 198
rect 113 168 145 198
rect 152 168 159 198
rect 66 116 71 146
rect 78 116 106 146
rect 113 136 121 146
rect 113 116 137 136
rect 35 50 37 80
rect 44 67 62 80
rect 44 50 50 67
rect 181 136 186 146
rect 165 116 186 136
rect 193 116 222 146
rect 229 136 234 146
rect 229 116 250 136
rect 88 67 106 80
rect 101 50 106 67
rect 113 50 145 80
rect 152 66 171 80
rect 327 168 333 198
rect 340 168 350 198
rect 290 116 292 146
rect 299 116 305 146
rect 152 50 155 66
rect 219 50 222 80
rect 229 50 260 80
rect 267 50 271 80
rect 66 8 71 38
rect 78 22 85 38
rect 78 8 101 22
rect 184 22 186 38
rect 168 8 186 22
rect 193 8 222 38
rect 229 8 233 38
<< pdiffusion >>
rect 65 448 71 496
rect 78 448 84 496
rect 100 448 106 496
rect 113 470 131 496
rect 113 448 115 470
rect 34 388 37 436
rect 44 409 62 436
rect 44 388 46 409
rect 219 448 222 496
rect 229 448 239 496
rect 255 448 260 496
rect 267 470 286 496
rect 267 448 270 470
rect 103 419 106 436
rect 87 388 106 419
rect 113 409 145 436
rect 113 388 117 409
rect 133 388 145 409
rect 152 388 165 436
rect 183 388 186 436
rect 193 404 222 436
rect 193 388 203 404
rect 219 388 222 404
rect 229 419 231 436
rect 229 388 242 419
rect 314 405 333 436
rect 330 388 333 405
rect 340 388 342 436
rect 49 326 71 352
rect 65 304 71 326
rect 78 304 87 352
rect 103 304 106 352
rect 113 304 116 352
rect 132 304 145 352
rect 152 304 165 352
rect 183 304 186 352
rect 193 326 222 352
rect 193 304 195 326
rect 211 304 222 326
rect 229 304 232 352
rect 289 304 292 352
rect 299 326 317 352
rect 299 304 301 326
<< ntransistor >>
rect 106 168 113 198
rect 145 168 152 198
rect 71 116 78 146
rect 106 116 113 146
rect 37 50 44 80
rect 186 116 193 146
rect 222 116 229 146
rect 106 50 113 80
rect 145 50 152 80
rect 333 168 340 198
rect 292 116 299 146
rect 222 50 229 80
rect 260 50 267 80
rect 71 8 78 38
rect 186 8 193 38
rect 222 8 229 38
<< ptransistor >>
rect 71 448 78 496
rect 106 448 113 496
rect 37 388 44 436
rect 222 448 229 496
rect 260 448 267 496
rect 106 388 113 436
rect 145 388 152 436
rect 186 388 193 436
rect 222 388 229 436
rect 333 388 340 436
rect 71 304 78 352
rect 106 304 113 352
rect 145 304 152 352
rect 186 304 193 352
rect 222 304 229 352
rect 292 304 299 352
<< polycontact >>
rect 98 579 123 604
rect 62 543 87 568
rect 29 506 54 531
rect 177 480 193 496
rect 177 446 193 462
rect 324 480 340 496
rect 283 388 299 404
rect 255 362 271 378
rect 140 278 156 294
rect 222 278 238 294
rect 222 90 238 106
rect 283 156 299 172
rect 177 50 193 66
rect 141 1 158 18
rect 260 8 276 39
rect 324 50 340 80
<< ndiffcontact >>
rect 88 168 104 198
rect 159 168 175 198
rect 50 116 66 146
rect 121 136 137 152
rect 19 50 35 80
rect 50 50 66 67
rect 165 136 181 152
rect 234 136 250 152
rect 85 50 101 67
rect 311 168 327 198
rect 350 168 366 198
rect 274 116 290 146
rect 305 116 321 146
rect 155 50 171 66
rect 203 50 219 80
rect 271 50 287 80
rect 50 8 66 38
rect 85 22 101 38
rect 168 22 184 38
rect 233 8 249 38
<< pdiffcontact >>
rect 49 448 65 496
rect 84 448 100 496
rect 115 448 131 470
rect 18 388 34 436
rect 46 388 62 409
rect 203 448 219 496
rect 239 448 255 496
rect 270 448 286 470
rect 87 419 103 436
rect 117 388 133 409
rect 165 388 183 436
rect 203 388 219 404
rect 231 419 247 436
rect 314 388 330 405
rect 342 388 358 436
rect 49 304 65 326
rect 87 304 103 352
rect 116 304 132 352
rect 165 304 183 352
rect 195 304 211 326
rect 232 304 248 352
rect 273 304 289 352
rect 301 304 317 326
<< psubstratetap >>
rect 118 212 136 228
<< nsubstratetap >>
rect 119 249 137 265
<< metal1 >>
rect 0 579 98 604
rect 123 579 372 604
rect 0 543 62 568
rect 87 543 372 568
rect 0 506 29 531
rect 54 506 372 531
rect 100 480 177 496
rect 49 436 65 448
rect 115 436 131 448
rect 34 419 87 436
rect 103 419 131 436
rect 141 446 177 462
rect 255 480 324 496
rect 141 409 154 446
rect 203 436 219 448
rect 270 436 286 448
rect 62 388 117 409
rect 133 388 154 409
rect 183 419 231 436
rect 247 419 342 436
rect 219 388 283 404
rect 18 352 34 388
rect 314 378 330 388
rect 116 362 255 378
rect 271 362 330 378
rect 116 352 132 362
rect 342 352 358 388
rect 18 336 87 352
rect 18 310 34 336
rect 19 268 34 310
rect 183 336 232 352
rect 248 336 273 352
rect 289 336 358 352
rect 49 294 65 304
rect 195 294 211 304
rect 301 294 317 304
rect 49 278 140 294
rect 156 278 211 294
rect 238 278 317 294
rect 342 268 358 336
rect 0 265 373 268
rect 0 249 119 265
rect 137 249 373 265
rect 0 243 373 249
rect 0 228 373 233
rect 0 212 118 228
rect 136 212 373 228
rect 0 208 373 212
rect 19 87 35 208
rect 88 198 104 208
rect 121 152 137 208
rect 175 182 311 198
rect 234 156 283 172
rect 234 152 250 156
rect 49 116 50 126
rect 137 136 165 152
rect 66 116 274 126
rect 305 106 321 116
rect 238 90 321 106
rect 19 80 219 87
rect 35 77 203 80
rect 66 50 85 67
rect 171 50 177 66
rect 287 50 324 80
rect 19 38 35 50
rect 350 39 366 168
rect 19 8 50 38
rect 101 28 168 38
rect 158 8 233 12
rect 276 8 366 39
rect 158 1 249 8
<< labels >>
rlabel metal1 373 243 373 268 7 Vdd!
rlabel metal1 373 208 373 233 7 GND!
rlabel metal1 0 243 0 268 3 Vdd!
rlabel metal1 0 208 0 233 3 GND!
rlabel metal1 372 579 372 604 7 nRst
rlabel metal1 372 543 372 568 7 Clk
rlabel metal1 372 506 372 531 7 D
rlabel metal1 0 579 0 604 3 nRst
rlabel metal1 0 543 0 568 3 Clk
rlabel metal1 0 506 0 531 3 D
rlabel polysilicon 333 610 340 610 5 Q
rlabel polysilicon 260 610 267 610 5 nQ
<< end >>
