magic
tech c035u
timestamp 1384420580
<< nwell >>
rect 0 124 111 220
<< polysilicon >>
rect 29 180 36 188
rect 56 180 63 188
rect 29 122 36 132
rect 56 122 63 132
rect 29 76 36 106
rect 56 76 63 106
rect 29 38 36 46
rect 56 38 63 46
<< ndiffusion >>
rect 27 46 29 76
rect 36 46 38 76
rect 54 46 56 76
rect 63 46 65 76
<< pdiffusion >>
rect 27 132 29 180
rect 36 132 56 180
rect 63 132 65 180
<< nohmic >>
rect 34 205 89 215
rect 34 199 68 205
<< ntransistor >>
rect 29 46 36 76
rect 56 46 63 76
<< ptransistor >>
rect 29 132 36 180
rect 56 132 63 180
<< polycontact >>
rect 22 106 38 122
rect 48 106 64 122
<< ndiffcontact >>
rect 3 46 27 76
rect 38 46 54 76
rect 65 46 89 76
<< pdiffcontact >>
rect 3 132 27 180
rect 65 132 91 180
<< nsubstratetap >>
rect 6 199 22 215
rect 89 199 105 215
<< metal1 >>
rect 0 199 6 215
rect 22 199 89 215
rect 105 199 111 215
rect 0 190 111 199
rect 3 180 27 190
rect 74 102 84 132
rect 44 86 74 96
rect 44 76 54 86
rect 3 36 27 46
rect 65 36 89 46
rect 3 10 111 36
<< m2contact >>
rect 74 86 90 102
<< metal2 >>
rect 24 0 36 220
rect 48 121 60 220
rect 48 0 60 107
rect 72 102 84 220
rect 72 86 74 102
rect 72 0 84 86
<< labels >>
rlabel metal2 24 0 36 0 1 A
rlabel metal2 24 220 36 220 5 A
rlabel metal1 0 190 0 215 3 Vdd!
rlabel metal1 111 11 111 36 7 GND!
rlabel metal1 111 190 111 215 7 Vdd!
rlabel metal2 48 220 60 220 5 B
rlabel metal2 48 0 60 0 1 B
rlabel metal2 72 0 84 0 1 Y
rlabel metal2 72 220 84 220 5 Y
<< end >>
