magic
tech c035u
timestamp 1385906574
<< nwell >>
rect 0 308 34 652
<< pohmic >>
rect 0 67 34 83
<< nohmic >>
rect 0 636 34 652
<< metal1 >>
rect 0 682 34 692
rect 0 662 34 672
rect 0 646 34 652
rect 0 632 10 646
rect 24 632 34 646
rect 0 627 34 632
rect 0 67 34 92
rect 0 47 34 57
rect 0 27 34 37
rect 0 7 34 17
<< m2contact >>
rect 10 632 24 646
<< metal2 >>
rect 11 646 23 699
rect 11 0 23 632
<< labels >>
rlabel metal1 34 67 34 92 7 GND!
rlabel metal1 34 47 34 57 7 Clock
rlabel metal1 34 27 34 37 7 Test
rlabel metal1 0 67 0 92 3 GND!
rlabel metal1 0 47 0 57 3 Clock
rlabel metal1 0 27 0 37 3 Test
rlabel metal2 11 0 23 0 1 Vdd!
rlabel metal1 0 7 0 17 3 nReset
rlabel metal1 34 7 34 17 7 nReset
rlabel metal1 34 627 34 652 7 Vdd!
rlabel metal1 0 627 0 652 3 Vdd!
rlabel metal1 34 682 34 692 7 ScanReturn
rlabel metal1 0 682 0 692 3 ScanReturn
rlabel metal2 11 699 23 699 5 Vdd!
rlabel metal1 0 662 0 672 3 Scan
rlabel metal1 34 662 34 672 7 Scan
<< end >>
