magic
tech c035u
timestamp 1385632638
<< metal1 >>
rect 11 792 21 809
rect 0 782 27 792
rect 0 759 27 769
rect 0 721 27 746
<< m2contact >>
rect 9 809 23 823
<< metal2 >>
rect 23 809 183 821
rect 51 799 63 809
rect 171 799 183 809
use inv inv_1
timestamp 1385631115
transform 1 0 27 0 1 0
box 0 0 120 799
use inv inv_0
timestamp 1385631115
transform 1 0 147 0 1 0
box 0 0 120 799
use rightend rightend_0
timestamp 1385632559
transform 1 0 267 0 1 0
box 0 0 292 799
<< labels >>
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 0 782 0 792 3 nScan
<< end >>
