magic
tech c035u
timestamp 1386087476
<< nwell >>
rect 0 401 744 799
<< pwell >>
rect 0 0 744 401
<< polysilicon >>
rect 240 681 245 697
rect 375 691 382 719
rect 405 691 412 719
rect 456 704 523 711
rect 52 671 59 679
rect 82 671 89 679
rect 112 671 119 679
rect 156 671 163 679
rect 186 671 193 679
rect 213 671 220 679
rect 240 671 247 681
rect 52 375 59 623
rect 82 553 89 623
rect 112 539 119 623
rect 156 553 163 623
rect 112 523 117 539
rect 82 381 89 505
rect 52 235 59 359
rect 82 335 89 365
rect 112 335 119 523
rect 156 381 163 505
rect 186 381 193 623
rect 213 501 220 623
rect 156 335 163 365
rect 112 319 117 335
rect 82 235 89 305
rect 112 235 119 319
rect 156 235 163 305
rect 186 235 193 365
rect 213 355 220 485
rect 213 235 220 339
rect 240 235 247 623
rect 342 610 349 621
rect 270 583 275 599
rect 270 553 277 583
rect 270 358 277 505
rect 342 388 349 562
rect 375 486 382 643
rect 405 612 412 643
rect 458 612 465 623
rect 499 612 506 645
rect 516 624 523 704
rect 561 691 568 719
rect 619 691 626 719
rect 561 624 568 643
rect 516 617 568 624
rect 561 612 568 617
rect 405 486 412 564
rect 458 486 465 564
rect 499 486 506 564
rect 561 486 568 564
rect 619 532 626 643
rect 687 612 694 675
rect 270 275 277 328
rect 275 259 277 275
rect 342 220 349 372
rect 375 331 382 438
rect 405 402 412 438
rect 458 428 465 438
rect 474 412 486 419
rect 405 395 446 402
rect 439 358 446 395
rect 479 358 486 412
rect 499 410 506 438
rect 561 428 568 438
rect 499 403 527 410
rect 520 358 527 403
rect 561 358 568 412
rect 375 288 382 315
rect 439 288 446 328
rect 52 197 59 205
rect 82 197 89 205
rect 112 197 119 205
rect 156 197 163 205
rect 186 197 193 205
rect 213 197 220 205
rect 240 197 247 205
rect 342 182 349 190
rect 375 161 382 258
rect 439 220 446 258
rect 479 220 486 328
rect 520 220 527 328
rect 561 255 568 328
rect 561 248 575 255
rect 561 225 575 232
rect 561 220 568 225
rect 619 220 626 516
rect 651 486 658 539
rect 651 358 658 438
rect 651 288 658 328
rect 375 110 382 131
rect 439 127 446 190
rect 479 128 486 190
rect 520 161 527 190
rect 561 161 568 190
rect 619 180 626 190
rect 619 142 626 150
rect 651 142 658 258
rect 687 227 694 564
rect 677 220 694 227
rect 684 190 691 195
rect 677 188 691 190
rect 684 180 691 188
rect 684 142 691 150
rect 520 120 527 131
rect 561 120 568 131
<< ndiffusion >>
rect 80 305 82 335
rect 89 305 91 335
rect 154 305 156 335
rect 163 305 165 335
rect 268 328 270 358
rect 277 328 279 358
rect 50 205 52 235
rect 59 205 82 235
rect 89 205 91 235
rect 107 205 112 235
rect 119 205 138 235
rect 154 205 156 235
rect 163 205 186 235
rect 193 205 195 235
rect 211 205 213 235
rect 220 205 240 235
rect 247 205 249 235
rect 434 328 439 358
rect 446 328 479 358
rect 486 328 493 358
rect 509 328 520 358
rect 527 328 561 358
rect 568 328 573 358
rect 370 258 375 288
rect 382 258 439 288
rect 446 258 457 288
rect 340 190 342 220
rect 349 190 354 220
rect 649 258 651 288
rect 658 258 664 288
rect 437 190 439 220
rect 446 190 479 220
rect 486 190 489 220
rect 553 190 561 220
rect 568 190 619 220
rect 626 190 630 220
rect 370 131 375 161
rect 382 131 387 161
rect 518 131 520 161
rect 527 131 561 161
rect 568 131 572 161
rect 681 150 684 180
rect 691 150 694 180
<< pdiffusion >>
rect 50 623 52 671
rect 59 623 64 671
rect 80 623 82 671
rect 89 623 91 671
rect 107 623 112 671
rect 119 623 138 671
rect 154 623 156 671
rect 163 623 165 671
rect 181 623 186 671
rect 193 623 195 671
rect 211 623 213 671
rect 220 623 222 671
rect 238 623 240 671
rect 247 623 249 671
rect 373 643 375 691
rect 382 643 384 691
rect 400 643 405 691
rect 412 643 414 691
rect 80 505 82 553
rect 89 505 91 553
rect 154 505 156 553
rect 163 505 165 553
rect 339 562 342 610
rect 349 562 354 610
rect 268 505 270 553
rect 277 505 279 553
rect 544 643 561 691
rect 568 643 578 691
rect 594 643 619 691
rect 626 643 629 691
rect 403 564 405 612
rect 412 564 440 612
rect 456 564 458 612
rect 465 564 475 612
rect 491 564 499 612
rect 506 564 508 612
rect 524 564 561 612
rect 568 564 570 612
rect 684 564 687 612
rect 694 564 704 612
rect 373 438 375 486
rect 382 438 385 486
rect 401 438 405 486
rect 412 438 414 486
rect 434 438 458 486
rect 465 438 473 486
rect 491 438 499 486
rect 506 438 508 486
rect 524 438 561 486
rect 568 438 571 486
rect 648 438 651 486
rect 658 438 664 486
<< pohmic >>
rect 0 79 30 86
rect 46 79 58 86
rect 74 79 86 86
rect 102 79 114 86
rect 130 79 142 86
rect 158 79 170 86
rect 186 79 198 86
rect 214 79 226 86
rect 242 79 254 86
rect 270 79 282 86
rect 298 79 318 86
rect 0 76 318 79
rect 334 76 346 86
rect 362 76 374 86
rect 390 76 402 86
rect 418 76 430 86
rect 446 76 458 86
rect 474 76 486 86
rect 502 76 514 86
rect 530 76 542 86
rect 559 76 571 86
rect 587 76 599 86
rect 615 76 627 86
rect 643 76 655 86
rect 672 76 684 86
rect 701 76 713 86
rect 730 76 744 86
<< nohmic >>
rect 0 743 318 746
rect 0 736 30 743
rect 46 736 58 743
rect 74 736 86 743
rect 102 736 114 743
rect 130 736 142 743
rect 158 736 170 743
rect 186 736 198 743
rect 214 736 226 743
rect 242 736 254 743
rect 270 736 282 743
rect 298 736 318 743
rect 334 736 346 746
rect 362 736 374 746
rect 390 736 402 746
rect 418 736 430 746
rect 446 736 458 746
rect 474 736 486 746
rect 502 736 514 746
rect 530 736 542 746
rect 558 736 570 746
rect 586 736 598 746
rect 614 736 626 746
rect 642 736 654 746
rect 670 736 682 746
rect 698 736 710 746
rect 726 736 744 746
<< ntransistor >>
rect 82 305 89 335
rect 156 305 163 335
rect 270 328 277 358
rect 52 205 59 235
rect 82 205 89 235
rect 112 205 119 235
rect 156 205 163 235
rect 186 205 193 235
rect 213 205 220 235
rect 240 205 247 235
rect 439 328 446 358
rect 479 328 486 358
rect 520 328 527 358
rect 561 328 568 358
rect 375 258 382 288
rect 439 258 446 288
rect 342 190 349 220
rect 651 258 658 288
rect 439 190 446 220
rect 479 190 486 220
rect 561 190 568 220
rect 619 190 626 220
rect 375 131 382 161
rect 520 131 527 161
rect 561 131 568 161
rect 684 150 691 180
<< ptransistor >>
rect 52 623 59 671
rect 82 623 89 671
rect 112 623 119 671
rect 156 623 163 671
rect 186 623 193 671
rect 213 623 220 671
rect 240 623 247 671
rect 375 643 382 691
rect 405 643 412 691
rect 82 505 89 553
rect 156 505 163 553
rect 342 562 349 610
rect 270 505 277 553
rect 561 643 568 691
rect 619 643 626 691
rect 405 564 412 612
rect 458 564 465 612
rect 499 564 506 612
rect 561 564 568 612
rect 687 564 694 612
rect 375 438 382 486
rect 405 438 412 486
rect 458 438 465 486
rect 499 438 506 486
rect 561 438 568 486
rect 651 438 658 486
<< polycontact >>
rect 245 681 261 697
rect 440 695 456 711
rect 490 645 506 661
rect 117 523 133 539
rect 48 359 64 375
rect 78 365 94 381
rect 204 485 220 501
rect 151 365 167 381
rect 182 365 198 381
rect 117 319 133 335
rect 204 339 220 355
rect 275 583 291 599
rect 678 675 694 691
rect 642 539 658 555
rect 614 516 630 532
rect 333 372 349 388
rect 259 259 275 275
rect 458 412 474 428
rect 561 412 577 428
rect 371 315 387 331
rect 563 232 579 248
rect 642 328 658 358
rect 511 190 527 220
rect 619 150 635 180
rect 668 190 684 220
rect 434 111 450 127
rect 475 111 492 128
<< ndiffcontact >>
rect 64 305 80 335
rect 91 305 107 335
rect 138 305 154 335
rect 165 305 181 335
rect 252 328 268 358
rect 279 328 295 358
rect 34 205 50 235
rect 91 205 107 235
rect 138 205 154 235
rect 195 205 211 235
rect 249 205 265 235
rect 418 328 434 358
rect 493 328 509 358
rect 573 328 589 358
rect 354 258 370 288
rect 457 258 473 288
rect 324 190 340 220
rect 354 190 370 220
rect 633 258 649 288
rect 664 258 680 288
rect 421 190 437 220
rect 489 190 505 220
rect 537 190 553 220
rect 630 190 646 220
rect 354 131 370 161
rect 387 131 403 161
rect 502 131 518 161
rect 572 131 588 161
rect 665 150 681 180
rect 694 150 710 180
<< pdiffcontact >>
rect 33 623 50 671
rect 64 623 80 671
rect 91 623 107 671
rect 138 623 154 671
rect 165 623 181 671
rect 195 623 211 671
rect 222 623 238 671
rect 249 623 265 671
rect 357 643 373 691
rect 384 643 400 691
rect 414 643 430 691
rect 64 505 80 553
rect 91 505 107 553
rect 138 505 154 553
rect 165 505 181 553
rect 323 562 339 610
rect 354 562 370 610
rect 252 505 268 553
rect 279 505 295 553
rect 528 643 544 691
rect 578 643 594 691
rect 629 643 645 691
rect 387 564 403 612
rect 440 564 456 612
rect 475 564 491 612
rect 508 564 524 612
rect 570 564 586 612
rect 668 564 684 612
rect 704 564 720 612
rect 357 438 373 486
rect 385 438 401 486
rect 414 438 434 486
rect 473 438 491 486
rect 508 438 524 486
rect 571 438 587 486
rect 632 438 648 486
rect 664 438 681 486
<< psubstratetap >>
rect 30 79 46 96
rect 58 79 74 96
rect 86 79 102 96
rect 114 79 130 96
rect 142 79 158 96
rect 170 79 186 96
rect 198 79 214 96
rect 226 79 242 96
rect 254 79 270 96
rect 282 79 298 96
rect 318 76 334 92
rect 346 76 362 92
rect 374 76 390 92
rect 402 76 418 92
rect 430 76 446 92
rect 458 76 474 92
rect 486 76 502 92
rect 514 76 530 92
rect 542 76 559 92
rect 571 76 587 92
rect 599 76 615 92
rect 627 76 643 92
rect 655 76 672 92
rect 684 76 701 92
rect 713 76 730 92
<< nsubstratetap >>
rect 30 727 46 743
rect 58 727 74 743
rect 86 727 102 743
rect 114 727 130 743
rect 142 727 158 743
rect 170 727 186 743
rect 198 727 214 743
rect 226 727 242 743
rect 254 727 270 743
rect 282 727 298 743
rect 318 730 334 746
rect 346 730 362 746
rect 374 730 390 746
rect 402 730 418 746
rect 430 730 446 746
rect 458 730 474 746
rect 486 730 502 746
rect 514 730 530 746
rect 542 730 558 746
rect 570 730 586 746
rect 598 730 614 746
rect 626 730 642 746
rect 654 730 670 746
rect 682 730 698 746
rect 710 730 726 746
<< metal1 >>
rect 0 782 744 792
rect 0 759 198 769
rect 276 759 622 769
rect 638 759 744 769
rect 0 743 318 746
rect 0 727 30 743
rect 46 727 58 743
rect 74 727 86 743
rect 102 727 114 743
rect 130 727 142 743
rect 158 727 170 743
rect 186 727 198 743
rect 214 727 226 743
rect 242 727 254 743
rect 270 727 282 743
rect 298 730 318 743
rect 334 730 346 746
rect 362 730 374 746
rect 390 730 402 746
rect 418 730 430 746
rect 446 730 458 746
rect 474 730 486 746
rect 502 730 514 746
rect 530 730 542 746
rect 558 730 570 746
rect 586 730 598 746
rect 614 730 626 746
rect 642 730 654 746
rect 670 730 682 746
rect 698 730 710 746
rect 726 730 744 746
rect 298 727 744 730
rect 0 721 744 727
rect 33 671 50 721
rect 91 671 107 721
rect 117 701 235 711
rect 39 573 50 623
rect 67 613 77 623
rect 117 613 127 701
rect 144 681 208 691
rect 144 671 154 681
rect 198 671 208 681
rect 225 671 235 701
rect 323 634 339 721
rect 357 691 373 721
rect 384 701 440 711
rect 384 691 400 701
rect 578 701 678 711
rect 578 691 594 701
rect 678 691 694 695
rect 323 633 340 634
rect 414 633 430 643
rect 67 603 127 613
rect 168 593 178 623
rect 198 613 208 623
rect 252 613 262 623
rect 198 603 262 613
rect 323 621 430 633
rect 440 645 490 655
rect 323 610 339 621
rect 387 612 403 621
rect 168 583 275 593
rect 39 563 262 573
rect 64 553 74 563
rect 169 553 181 563
rect 133 523 138 539
rect 252 553 262 563
rect 97 495 107 505
rect 97 485 204 495
rect 285 385 295 505
rect 323 511 339 562
rect 440 612 456 645
rect 528 633 544 643
rect 629 633 645 643
rect 704 633 720 721
rect 475 623 720 633
rect 475 612 491 623
rect 570 612 586 623
rect 704 612 720 623
rect 354 549 370 562
rect 440 549 456 564
rect 354 539 456 549
rect 508 554 524 564
rect 508 544 642 554
rect 414 516 574 526
rect 590 516 614 526
rect 668 526 684 564
rect 630 516 684 526
rect 323 501 401 511
rect 385 486 401 501
rect 414 486 434 516
rect 704 506 720 564
rect 473 496 587 506
rect 473 486 491 496
rect 571 486 587 496
rect 632 496 720 506
rect 632 486 648 496
rect 587 438 632 486
rect 357 428 373 438
rect 508 428 524 438
rect 664 428 681 438
rect 357 418 458 428
rect 474 418 524 428
rect 577 418 681 428
rect 372 390 509 402
rect 144 365 151 379
rect 285 375 333 385
rect 285 358 295 375
rect 97 345 204 355
rect 97 335 107 345
rect 133 319 138 335
rect 70 295 80 305
rect 171 295 181 305
rect 372 353 385 390
rect 493 358 509 390
rect 324 341 385 353
rect 252 295 262 328
rect 70 285 295 295
rect 37 265 259 275
rect 37 235 47 265
rect 94 245 174 255
rect 94 235 104 245
rect 138 101 154 205
rect 164 195 174 245
rect 198 235 208 265
rect 252 195 262 205
rect 164 185 262 195
rect 285 101 295 285
rect 324 288 340 341
rect 371 314 387 315
rect 589 328 642 358
rect 418 318 434 328
rect 418 308 710 318
rect 324 258 354 288
rect 473 278 633 288
rect 324 220 340 258
rect 354 247 370 258
rect 664 248 680 258
rect 354 235 553 247
rect 537 220 553 235
rect 579 232 680 248
rect 370 190 421 220
rect 505 190 511 220
rect 646 190 668 220
rect 324 161 340 190
rect 694 180 710 308
rect 324 131 354 161
rect 403 151 502 161
rect 635 150 665 180
rect 324 101 342 131
rect 433 111 434 127
rect 572 121 588 131
rect 492 111 588 121
rect 0 96 744 101
rect 0 79 30 96
rect 46 79 58 96
rect 74 79 86 96
rect 102 79 114 96
rect 130 79 142 96
rect 158 79 170 96
rect 186 79 198 96
rect 214 79 226 96
rect 242 79 254 96
rect 270 79 282 96
rect 298 92 744 96
rect 298 79 318 92
rect 0 76 318 79
rect 334 76 346 92
rect 362 76 374 92
rect 390 76 402 92
rect 418 76 430 92
rect 446 76 458 92
rect 474 76 486 92
rect 502 76 514 92
rect 530 76 542 92
rect 559 76 571 92
rect 587 76 599 92
rect 615 76 627 92
rect 643 76 655 92
rect 672 76 684 92
rect 701 76 713 92
rect 730 76 744 92
rect 0 53 371 63
rect 387 53 744 63
rect 0 30 130 40
rect 144 30 744 40
rect 0 7 417 17
rect 433 7 744 17
<< m2contact >>
rect 198 757 212 771
rect 262 758 276 772
rect 622 756 638 772
rect 261 683 275 697
rect 678 695 694 711
rect 574 516 590 532
rect 94 367 109 381
rect 130 365 144 379
rect 198 367 212 381
rect 48 345 62 359
rect 371 298 387 314
rect 417 111 433 127
rect 371 50 387 66
rect 130 28 144 42
rect 417 3 433 19
<< metal2 >>
rect 48 359 60 799
rect 96 381 108 799
rect 199 743 211 757
rect 198 727 211 743
rect 199 381 211 727
rect 263 697 275 758
rect 576 532 588 799
rect 624 772 636 799
rect 624 711 636 756
rect 624 695 678 711
rect 48 0 60 345
rect 96 0 108 367
rect 131 42 143 365
rect 371 66 387 298
rect 417 19 433 111
rect 576 0 588 516
rect 624 0 636 695
<< labels >>
rlabel metal2 48 799 60 799 5 D
rlabel metal2 48 0 60 0 1 D
rlabel metal2 96 0 108 0 1 Load
rlabel metal2 96 799 108 799 5 Load
rlabel metal2 576 799 588 799 5 nQ
rlabel metal2 576 0 588 0 1 nQ
rlabel metal2 624 799 636 799 5 Q
rlabel metal2 624 0 636 0 1 Q
rlabel metal1 744 782 744 792 7 ScanReturn
rlabel metal1 744 759 744 769 7 Q
rlabel metal1 744 76 744 101 7 GND!
rlabel metal1 744 53 744 63 7 Clock
rlabel metal1 744 30 744 40 7 Test
rlabel metal1 744 7 744 17 7 nReset
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 53 0 63 3 Clock
<< end >>
