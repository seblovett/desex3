magic
tech c035u
timestamp 1384960332
<< nwell >>
rect 0 517 144 729
<< metal1 >>
rect 0 765 144 775
rect 0 742 144 752
rect 0 704 144 729
rect 0 69 144 94
rect 0 46 144 56
rect 0 23 144 33
rect 0 0 144 10
<< labels >>
rlabel metal1 0 0 0 10 2 nReset
rlabel metal1 144 0 144 10 8 nReset
rlabel metal1 0 23 0 33 3 Test
rlabel metal1 144 23 144 33 7 Test
rlabel metal1 0 46 0 56 3 Clock
rlabel metal1 144 46 144 56 7 Clock
rlabel metal1 144 69 144 94 7 GND!
rlabel metal1 0 69 0 94 3 GND!
rlabel metal1 144 704 144 729 7 Vdd!
rlabel metal1 0 704 0 729 3 Vdd!
rlabel metal1 144 742 144 752 7 Scan
rlabel metal1 0 742 0 752 3 Scan
rlabel metal1 0 765 0 775 4 ScanReturn
rlabel metal1 144 765 144 775 6 ScanReturn
<< end >>
