magic
tech c035u
timestamp 1386264609
<< nwell >>
rect 20 445 1292 843
<< pwell >>
rect 20 44 1292 445
<< polysilicon >>
rect 87 735 94 763
rect 117 735 124 763
rect 168 748 235 755
rect 54 654 61 665
rect 54 432 61 606
rect 87 530 94 687
rect 117 656 124 687
rect 170 656 177 667
rect 211 656 218 689
rect 228 668 235 748
rect 273 735 280 763
rect 331 735 338 763
rect 273 668 280 687
rect 228 661 280 668
rect 273 656 280 661
rect 117 530 124 608
rect 170 530 177 608
rect 211 530 218 608
rect 273 530 280 608
rect 331 576 338 687
rect 399 656 406 719
rect 54 269 61 416
rect 87 375 94 482
rect 117 446 124 482
rect 170 472 177 482
rect 186 456 198 463
rect 117 439 158 446
rect 151 402 158 439
rect 191 402 198 456
rect 211 454 218 482
rect 273 472 280 482
rect 211 447 239 454
rect 232 402 239 447
rect 273 402 280 456
rect 87 332 94 359
rect 151 332 158 372
rect 54 231 61 239
rect 87 205 94 302
rect 151 269 158 302
rect 191 269 198 372
rect 232 269 239 372
rect 273 299 280 372
rect 273 292 287 299
rect 273 269 287 276
rect 273 264 280 269
rect 331 264 338 560
rect 363 530 370 583
rect 363 402 370 482
rect 363 332 370 372
rect 87 154 94 175
rect 151 171 158 239
rect 191 172 198 239
rect 232 205 239 239
rect 273 205 280 234
rect 331 224 338 234
rect 331 186 338 194
rect 363 186 370 302
rect 399 271 406 608
rect 507 513 514 521
rect 627 513 634 521
rect 747 513 754 521
rect 867 513 874 521
rect 987 513 994 521
rect 1107 513 1114 521
rect 1227 513 1234 521
rect 507 435 514 465
rect 627 435 634 465
rect 747 435 754 465
rect 867 435 874 465
rect 987 435 994 465
rect 1107 435 1114 465
rect 1227 435 1234 465
rect 512 419 514 435
rect 632 419 634 435
rect 752 419 754 435
rect 872 419 874 435
rect 992 419 994 435
rect 1112 419 1114 435
rect 1232 419 1234 435
rect 507 384 514 419
rect 627 384 634 419
rect 747 384 754 419
rect 867 384 874 419
rect 987 384 994 419
rect 1107 384 1114 419
rect 1227 384 1234 419
rect 507 346 514 354
rect 627 346 634 354
rect 747 346 754 354
rect 867 346 874 354
rect 987 346 994 354
rect 1107 346 1114 354
rect 1227 346 1234 354
rect 389 264 406 271
rect 396 234 403 239
rect 389 232 403 234
rect 396 224 403 232
rect 396 186 403 194
rect 232 164 239 175
rect 273 164 280 175
<< ndiffusion >>
rect 146 372 151 402
rect 158 372 191 402
rect 198 372 205 402
rect 221 372 232 402
rect 239 372 273 402
rect 280 372 285 402
rect 82 302 87 332
rect 94 302 151 332
rect 158 302 169 332
rect 52 239 54 269
rect 61 239 66 269
rect 149 239 151 269
rect 158 239 191 269
rect 198 239 201 269
rect 361 302 363 332
rect 370 302 376 332
rect 82 175 87 205
rect 94 175 99 205
rect 265 234 273 264
rect 280 234 331 264
rect 338 234 342 264
rect 230 175 232 205
rect 239 175 273 205
rect 280 175 284 205
rect 505 354 507 384
rect 514 354 516 384
rect 625 354 627 384
rect 634 354 636 384
rect 745 354 747 384
rect 754 354 756 384
rect 865 354 867 384
rect 874 354 876 384
rect 985 354 987 384
rect 994 354 996 384
rect 1105 354 1107 384
rect 1114 354 1116 384
rect 1225 354 1227 384
rect 1234 354 1236 384
rect 393 194 396 224
rect 403 194 406 224
<< pdiffusion >>
rect 85 687 87 735
rect 94 687 96 735
rect 112 687 117 735
rect 124 687 126 735
rect 51 606 54 654
rect 61 606 66 654
rect 256 687 273 735
rect 280 687 290 735
rect 306 687 331 735
rect 338 687 341 735
rect 115 608 117 656
rect 124 608 152 656
rect 168 608 170 656
rect 177 608 187 656
rect 203 608 211 656
rect 218 608 220 656
rect 236 608 273 656
rect 280 608 282 656
rect 396 608 399 656
rect 406 608 416 656
rect 85 482 87 530
rect 94 482 97 530
rect 113 482 117 530
rect 124 482 126 530
rect 146 482 170 530
rect 177 482 185 530
rect 203 482 211 530
rect 218 482 220 530
rect 236 482 273 530
rect 280 482 283 530
rect 360 482 363 530
rect 370 482 376 530
rect 505 465 507 513
rect 514 465 516 513
rect 625 465 627 513
rect 634 465 636 513
rect 745 465 747 513
rect 754 465 756 513
rect 865 465 867 513
rect 874 465 876 513
rect 985 465 987 513
rect 994 465 996 513
rect 1105 465 1107 513
rect 1114 465 1116 513
rect 1225 465 1227 513
rect 1234 465 1236 513
<< pohmic >>
rect 20 120 30 130
rect 46 120 58 130
rect 74 120 86 130
rect 102 120 114 130
rect 130 120 142 130
rect 158 120 170 130
rect 186 120 198 130
rect 214 120 226 130
rect 242 120 254 130
rect 271 120 283 130
rect 299 120 311 130
rect 327 120 339 130
rect 355 120 367 130
rect 384 120 396 130
rect 413 120 425 130
rect 442 120 458 130
rect 474 120 486 130
rect 502 120 514 130
rect 530 120 542 130
rect 558 120 578 130
rect 594 120 606 130
rect 622 120 634 130
rect 650 120 662 130
rect 678 120 698 130
rect 714 120 726 130
rect 742 120 754 130
rect 770 120 782 130
rect 798 120 818 130
rect 834 120 846 130
rect 862 120 874 130
rect 890 120 902 130
rect 918 120 938 130
rect 954 120 966 130
rect 982 120 994 130
rect 1010 120 1022 130
rect 1038 120 1058 130
rect 1074 120 1086 130
rect 1102 120 1114 130
rect 1130 120 1142 130
rect 1158 120 1178 130
rect 1194 120 1206 130
rect 1222 120 1234 130
rect 1250 120 1262 130
rect 1278 120 1292 130
<< nohmic >>
rect 20 780 30 790
rect 46 780 58 790
rect 74 780 86 790
rect 102 780 114 790
rect 130 780 142 790
rect 158 780 170 790
rect 186 780 198 790
rect 214 780 226 790
rect 242 780 254 790
rect 270 780 282 790
rect 298 780 310 790
rect 326 780 338 790
rect 354 780 366 790
rect 382 780 394 790
rect 410 780 422 790
rect 438 780 458 790
rect 474 780 486 790
rect 502 780 514 790
rect 530 780 542 790
rect 558 780 578 790
rect 594 780 606 790
rect 622 780 634 790
rect 650 780 662 790
rect 678 780 698 790
rect 714 780 726 790
rect 742 780 754 790
rect 770 780 782 790
rect 798 780 818 790
rect 834 780 846 790
rect 862 780 874 790
rect 890 780 902 790
rect 918 780 938 790
rect 954 780 966 790
rect 982 780 994 790
rect 1010 780 1022 790
rect 1038 780 1058 790
rect 1074 780 1086 790
rect 1102 780 1114 790
rect 1130 780 1142 790
rect 1158 780 1178 790
rect 1194 780 1206 790
rect 1222 780 1234 790
rect 1250 780 1262 790
rect 1278 780 1292 790
<< ntransistor >>
rect 151 372 158 402
rect 191 372 198 402
rect 232 372 239 402
rect 273 372 280 402
rect 87 302 94 332
rect 151 302 158 332
rect 54 239 61 269
rect 151 239 158 269
rect 191 239 198 269
rect 363 302 370 332
rect 87 175 94 205
rect 273 234 280 264
rect 331 234 338 264
rect 232 175 239 205
rect 273 175 280 205
rect 507 354 514 384
rect 627 354 634 384
rect 747 354 754 384
rect 867 354 874 384
rect 987 354 994 384
rect 1107 354 1114 384
rect 1227 354 1234 384
rect 396 194 403 224
<< ptransistor >>
rect 87 687 94 735
rect 117 687 124 735
rect 54 606 61 654
rect 273 687 280 735
rect 331 687 338 735
rect 117 608 124 656
rect 170 608 177 656
rect 211 608 218 656
rect 273 608 280 656
rect 399 608 406 656
rect 87 482 94 530
rect 117 482 124 530
rect 170 482 177 530
rect 211 482 218 530
rect 273 482 280 530
rect 363 482 370 530
rect 507 465 514 513
rect 627 465 634 513
rect 747 465 754 513
rect 867 465 874 513
rect 987 465 994 513
rect 1107 465 1114 513
rect 1227 465 1234 513
<< polycontact >>
rect 152 739 168 755
rect 202 689 218 705
rect 390 719 406 735
rect 354 583 370 599
rect 326 560 342 576
rect 45 416 61 432
rect 170 456 186 472
rect 273 456 289 472
rect 83 359 99 375
rect 275 276 291 292
rect 223 239 239 269
rect 354 372 370 402
rect 331 194 347 224
rect 496 419 512 435
rect 616 419 632 435
rect 736 419 752 435
rect 856 419 872 435
rect 976 419 992 435
rect 1096 419 1112 435
rect 1216 419 1232 435
rect 380 234 396 264
rect 146 155 162 171
rect 187 155 204 172
<< ndiffcontact >>
rect 130 372 146 402
rect 205 372 221 402
rect 285 372 301 402
rect 66 302 82 332
rect 169 302 185 332
rect 36 239 52 269
rect 66 239 82 269
rect 133 239 149 269
rect 201 239 217 269
rect 345 302 361 332
rect 376 302 392 332
rect 66 175 82 205
rect 99 175 115 205
rect 249 234 265 264
rect 342 234 358 264
rect 214 175 230 205
rect 284 175 300 205
rect 489 354 505 384
rect 516 354 532 384
rect 609 354 625 384
rect 636 354 652 384
rect 729 354 745 384
rect 756 354 772 384
rect 849 354 865 384
rect 876 354 892 384
rect 969 354 985 384
rect 996 354 1012 384
rect 1089 354 1105 384
rect 1116 354 1132 384
rect 1209 354 1225 384
rect 1236 354 1252 384
rect 377 194 393 224
rect 406 194 422 224
<< pdiffcontact >>
rect 69 687 85 735
rect 96 687 112 735
rect 126 687 142 735
rect 35 606 51 654
rect 66 606 82 654
rect 240 687 256 735
rect 290 687 306 735
rect 341 687 357 735
rect 99 608 115 656
rect 152 608 168 656
rect 187 608 203 656
rect 220 608 236 656
rect 282 608 298 656
rect 380 608 396 656
rect 416 608 432 656
rect 69 482 85 530
rect 97 482 113 530
rect 126 482 146 530
rect 185 482 203 530
rect 220 482 236 530
rect 283 482 299 530
rect 344 482 360 530
rect 376 482 393 530
rect 489 465 505 513
rect 516 465 532 513
rect 609 465 625 513
rect 636 465 652 513
rect 729 465 745 513
rect 756 465 772 513
rect 849 465 865 513
rect 876 465 892 513
rect 969 465 985 513
rect 996 465 1012 513
rect 1089 465 1105 513
rect 1116 465 1132 513
rect 1209 465 1225 513
rect 1236 465 1252 513
<< psubstratetap >>
rect 33 381 49 397
rect 36 210 52 226
rect 489 325 505 341
rect 609 325 625 341
rect 729 325 745 341
rect 849 325 865 341
rect 969 325 985 341
rect 1089 325 1105 341
rect 1209 325 1225 341
rect 30 120 46 136
rect 58 120 74 136
rect 86 120 102 136
rect 114 120 130 136
rect 142 120 158 136
rect 170 120 186 136
rect 198 120 214 136
rect 226 120 242 136
rect 254 120 271 136
rect 283 120 299 136
rect 311 120 327 136
rect 339 120 355 136
rect 367 120 384 136
rect 396 120 413 136
rect 425 120 442 136
rect 458 120 474 136
rect 486 120 502 136
rect 514 120 530 136
rect 542 120 558 136
rect 578 120 594 136
rect 606 120 622 136
rect 634 120 650 136
rect 662 120 678 136
rect 698 120 714 136
rect 726 120 742 136
rect 754 120 770 136
rect 782 120 798 136
rect 818 120 834 136
rect 846 120 862 136
rect 874 120 890 136
rect 902 120 918 136
rect 938 120 954 136
rect 966 120 982 136
rect 994 120 1010 136
rect 1022 120 1038 136
rect 1058 120 1074 136
rect 1086 120 1102 136
rect 1114 120 1130 136
rect 1142 120 1158 136
rect 1178 120 1194 136
rect 1206 120 1222 136
rect 1234 120 1250 136
rect 1262 120 1278 136
<< nsubstratetap >>
rect 30 774 46 790
rect 58 774 74 790
rect 86 774 102 790
rect 114 774 130 790
rect 142 774 158 790
rect 170 774 186 790
rect 198 774 214 790
rect 226 774 242 790
rect 254 774 270 790
rect 282 774 298 790
rect 310 774 326 790
rect 338 774 354 790
rect 366 774 382 790
rect 394 774 410 790
rect 422 774 438 790
rect 458 774 474 790
rect 486 774 502 790
rect 514 774 530 790
rect 542 774 558 790
rect 578 774 594 790
rect 606 774 622 790
rect 634 774 650 790
rect 662 774 678 790
rect 698 774 714 790
rect 726 774 742 790
rect 754 774 770 790
rect 782 774 798 790
rect 818 774 834 790
rect 846 774 862 790
rect 874 774 890 790
rect 902 774 918 790
rect 938 774 954 790
rect 966 774 982 790
rect 994 774 1010 790
rect 1022 774 1038 790
rect 1058 774 1074 790
rect 1086 774 1102 790
rect 1114 774 1130 790
rect 1142 774 1158 790
rect 1178 774 1194 790
rect 1206 774 1222 790
rect 1234 774 1250 790
rect 1262 774 1278 790
<< metal1 >>
rect 0 903 1003 914
rect 0 429 10 903
rect 298 875 714 885
rect 731 875 834 885
rect 347 851 474 861
rect 491 851 593 861
rect 20 826 1292 836
rect 20 803 330 813
rect 346 803 1292 813
rect 20 774 30 790
rect 46 774 58 790
rect 74 774 86 790
rect 102 774 114 790
rect 130 774 142 790
rect 158 774 170 790
rect 186 774 198 790
rect 214 774 226 790
rect 242 774 254 790
rect 270 774 282 790
rect 298 774 310 790
rect 326 774 338 790
rect 354 774 366 790
rect 382 774 394 790
rect 410 774 422 790
rect 438 774 458 790
rect 474 774 486 790
rect 502 774 514 790
rect 530 774 542 790
rect 558 774 578 790
rect 594 774 606 790
rect 622 774 634 790
rect 650 774 662 790
rect 678 774 698 790
rect 714 774 726 790
rect 742 774 754 790
rect 770 774 782 790
rect 798 774 818 790
rect 834 774 846 790
rect 862 774 874 790
rect 890 774 902 790
rect 918 774 938 790
rect 954 774 966 790
rect 982 774 994 790
rect 1010 774 1022 790
rect 1038 774 1058 790
rect 1074 774 1086 790
rect 1102 774 1114 790
rect 1130 774 1142 790
rect 1158 774 1178 790
rect 1194 774 1206 790
rect 1222 774 1234 790
rect 1250 774 1262 790
rect 1278 774 1328 790
rect 20 765 1328 774
rect 35 678 51 765
rect 69 735 85 765
rect 96 745 152 755
rect 96 735 112 745
rect 290 745 390 755
rect 290 735 306 745
rect 390 735 406 739
rect 35 677 52 678
rect 126 677 142 687
rect 35 665 142 677
rect 152 689 202 699
rect 35 654 51 665
rect 99 656 115 665
rect 35 555 51 606
rect 152 656 168 689
rect 240 677 256 687
rect 341 677 357 687
rect 416 677 432 765
rect 187 667 432 677
rect 187 656 203 667
rect 282 656 298 667
rect 416 656 432 667
rect 66 593 82 606
rect 152 593 168 608
rect 66 583 168 593
rect 220 598 236 608
rect 220 588 354 598
rect 126 560 282 570
rect 298 560 326 570
rect 380 570 396 608
rect 342 560 396 570
rect 35 545 113 555
rect 97 530 113 545
rect 126 530 146 560
rect 416 550 432 608
rect 185 540 299 550
rect 185 530 203 540
rect 283 530 299 540
rect 344 540 432 550
rect 344 530 360 540
rect 299 482 344 530
rect 69 472 85 482
rect 220 472 236 482
rect 376 472 393 482
rect 69 462 170 472
rect 186 462 236 472
rect 289 462 393 472
rect 489 513 505 765
rect 609 513 625 765
rect 729 513 745 765
rect 849 513 865 765
rect 969 513 985 765
rect 1089 513 1105 765
rect 1209 513 1225 765
rect 84 434 221 446
rect 0 419 45 429
rect 84 397 97 434
rect 205 402 221 434
rect 522 433 532 465
rect 642 433 652 465
rect 762 433 772 465
rect 882 433 892 465
rect 1002 433 1012 465
rect 1122 433 1132 465
rect 1242 433 1252 465
rect 49 385 97 397
rect 49 381 52 385
rect 36 332 52 381
rect 83 358 99 359
rect 301 372 354 402
rect 522 384 532 419
rect 642 384 652 419
rect 762 384 772 419
rect 882 384 892 419
rect 1002 384 1012 419
rect 1122 384 1132 419
rect 1242 384 1252 419
rect 130 362 146 372
rect 130 352 422 362
rect 36 302 66 332
rect 185 322 345 332
rect 36 269 52 302
rect 66 291 82 302
rect 376 292 392 302
rect 66 279 265 291
rect 82 239 133 269
rect 217 239 223 269
rect 249 264 265 279
rect 291 276 392 292
rect 36 226 52 239
rect 358 234 380 264
rect 406 224 422 352
rect 36 205 52 210
rect 36 175 66 205
rect 115 195 214 205
rect 347 194 377 224
rect 489 341 505 354
rect 36 145 54 175
rect 145 155 146 171
rect 284 165 300 175
rect 204 155 300 165
rect 489 145 505 325
rect 609 341 625 354
rect 609 145 625 325
rect 729 341 745 354
rect 729 145 745 325
rect 849 341 865 354
rect 849 145 865 325
rect 969 341 985 354
rect 969 145 985 325
rect 1089 341 1105 354
rect 1089 145 1105 325
rect 1209 341 1225 354
rect 1209 145 1225 325
rect 20 136 1328 145
rect 20 120 30 136
rect 46 120 58 136
rect 74 120 86 136
rect 102 120 114 136
rect 130 120 142 136
rect 158 120 170 136
rect 186 120 198 136
rect 214 120 226 136
rect 242 120 254 136
rect 271 120 283 136
rect 299 120 311 136
rect 327 120 339 136
rect 355 120 367 136
rect 384 120 396 136
rect 413 120 425 136
rect 442 120 458 136
rect 474 120 486 136
rect 502 120 514 136
rect 530 120 542 136
rect 558 120 578 136
rect 594 120 606 136
rect 622 120 634 136
rect 650 120 662 136
rect 678 120 698 136
rect 714 120 726 136
rect 742 120 754 136
rect 770 120 782 136
rect 798 120 818 136
rect 834 120 846 136
rect 862 120 874 136
rect 890 120 902 136
rect 918 120 938 136
rect 954 120 966 136
rect 982 120 994 136
rect 1010 120 1022 136
rect 1038 120 1058 136
rect 1074 120 1086 136
rect 1102 120 1114 136
rect 1130 120 1142 136
rect 1158 120 1178 136
rect 1194 120 1206 136
rect 1222 120 1234 136
rect 1250 120 1262 136
rect 1278 120 1328 136
rect 20 97 83 107
rect 99 97 1328 107
rect 20 74 1292 84
rect 20 51 129 61
rect 145 51 1308 61
rect 1298 34 1308 51
rect 1257 24 1308 34
rect 1318 12 1328 97
rect 1137 2 1328 12
<< m2contact >>
rect 1003 901 1017 915
rect 281 872 298 888
rect 714 872 731 888
rect 834 872 851 888
rect 330 850 347 864
rect 474 849 491 865
rect 593 849 610 865
rect 330 800 346 816
rect 390 739 406 755
rect 282 560 298 576
rect 482 420 496 434
rect 522 419 536 433
rect 602 420 616 434
rect 642 419 656 433
rect 722 420 736 434
rect 762 419 776 433
rect 842 420 856 434
rect 882 419 896 433
rect 962 420 976 434
rect 1002 419 1016 433
rect 1082 420 1096 434
rect 1122 419 1136 433
rect 1202 420 1216 434
rect 1242 419 1256 433
rect 83 342 99 358
rect 129 155 145 171
rect 83 94 99 110
rect 129 48 145 64
rect 1243 22 1257 36
rect 1123 0 1137 14
<< metal2 >>
rect 284 888 296 941
rect 284 576 296 872
rect 332 864 344 941
rect 332 816 344 850
rect 332 755 344 800
rect 332 739 390 755
rect 83 110 99 342
rect 129 64 145 155
rect 284 44 296 560
rect 332 44 344 739
rect 476 434 488 849
rect 476 420 482 434
rect 524 433 536 843
rect 476 44 488 420
rect 524 44 536 419
rect 596 434 608 849
rect 596 420 602 434
rect 644 433 656 843
rect 596 44 608 420
rect 644 44 656 419
rect 716 434 728 872
rect 716 420 722 434
rect 764 433 776 843
rect 716 44 728 420
rect 764 44 776 419
rect 836 434 848 872
rect 836 420 842 434
rect 884 433 896 843
rect 836 44 848 420
rect 884 44 896 419
rect 956 434 968 941
rect 1004 915 1016 941
rect 956 420 962 434
rect 1004 433 1016 901
rect 956 44 968 420
rect 1004 44 1016 419
rect 1076 434 1088 941
rect 1076 420 1082 434
rect 1124 433 1136 941
rect 1076 44 1088 420
rect 1124 14 1136 419
rect 1196 434 1208 941
rect 1196 420 1202 434
rect 1244 433 1256 941
rect 1196 44 1208 420
rect 1244 36 1256 419
<< labels >>
rlabel metal2 956 941 968 941 5 nD
rlabel metal2 284 941 296 941 5 nQ
rlabel metal2 332 941 344 941 5 Q
rlabel metal2 1196 941 1208 941 5 nnReset
rlabel metal2 1076 941 1088 941 5 nClock
rlabel metal1 1328 765 1328 790 7 Vdd!
rlabel metal1 1328 120 1328 145 7 GND!
rlabel metal2 1124 941 1136 941 1 Clock
rlabel metal2 1004 941 1016 941 5 D
rlabel metal2 1244 941 1256 941 5 nReset
<< end >>
