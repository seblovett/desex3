magic
tech c035u
timestamp 1386278660
<< pwell >>
rect 1824 159 1858 184
<< metal1 >>
rect 229 900 2669 910
rect 2683 900 2790 910
rect 2971 905 3035 915
rect 3025 875 3035 905
rect 1824 865 1858 875
rect 2098 865 2132 875
rect 2372 865 2406 875
rect 3006 865 3068 875
rect 1824 842 1858 852
rect 2098 842 2132 852
rect 2372 842 2406 852
rect 1824 804 1858 829
rect 2098 804 2132 829
rect 2372 804 2406 829
rect 1824 159 1858 184
rect 2098 159 2132 184
rect 2372 159 2406 184
rect 3006 159 3068 184
rect 1824 136 1833 146
rect 1847 136 1858 146
rect 2098 136 2132 146
rect 2372 136 2406 146
rect 3006 136 3068 146
rect 1824 113 1858 123
rect 2098 113 2108 123
rect 2122 113 2132 123
rect 2372 113 2406 123
rect 3006 113 3068 123
rect 1824 90 1858 100
rect 2098 90 2132 100
rect 2372 90 2381 100
rect 2395 90 2406 100
rect 3006 90 3068 100
rect 253 57 1535 67
rect 277 35 1655 45
rect 301 13 1775 23
<< m2contact >>
rect 215 898 229 912
rect 2669 898 2683 912
rect 2790 898 2804 912
rect 2957 901 2971 915
rect 1833 134 1847 148
rect 2108 111 2122 125
rect 2381 88 2395 102
rect 239 55 253 69
rect 1535 57 1549 71
rect 263 33 277 47
rect 1655 33 1669 47
rect 287 11 301 25
rect 1775 11 1789 25
<< metal2 >>
rect 216 912 228 945
rect 216 882 228 898
rect 2670 882 2682 898
rect 2790 882 2802 898
rect 2958 882 2970 901
rect 0 0 200 83
rect 216 0 228 83
rect 240 69 252 83
rect 240 0 252 55
rect 264 47 276 83
rect 264 0 276 33
rect 288 25 300 83
rect 288 0 300 11
rect 1488 0 1500 83
rect 1536 71 1548 83
rect 1608 0 1620 83
rect 1656 47 1668 83
rect 1728 0 1740 83
rect 1776 25 1788 83
rect 1835 71 1847 134
rect 1882 71 1894 83
rect 2002 71 2014 83
rect 1835 59 2014 71
rect 2108 72 2120 111
rect 2156 72 2168 83
rect 2276 72 2288 83
rect 2108 60 2288 72
rect 2383 73 2395 88
rect 2430 73 2442 83
rect 2550 73 2562 83
rect 2383 61 2562 73
rect 2910 0 2922 83
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 0 0 1 83
box 0 0 1464 799
use inv inv_0
timestamp 1386238110
transform 1 0 1464 0 1 83
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 1584 0 1 83
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 1704 0 1 83
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 1858 0 1 83
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 1978 0 1 83
box 0 0 120 799
use inv inv_5
timestamp 1386238110
transform 1 0 2132 0 1 83
box 0 0 120 799
use inv inv_6
timestamp 1386238110
transform 1 0 2252 0 1 83
box 0 0 120 799
use inv inv_7
timestamp 1386238110
transform 1 0 2406 0 1 83
box 0 0 120 799
use inv inv_8
timestamp 1386238110
transform 1 0 2526 0 1 83
box 0 0 120 799
use inv inv_9
timestamp 1386238110
transform 1 0 2646 0 1 83
box 0 0 120 799
use inv inv_10
timestamp 1386238110
transform 1 0 2766 0 1 83
box 0 0 120 799
use inv inv_11
timestamp 1386238110
transform 1 0 2886 0 1 83
box 0 0 120 799
<< labels >>
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 1488 0 1500 0 1 nTest
rlabel metal2 1608 0 1620 0 1 nClock
rlabel metal2 1728 0 1740 0 1 nnReset
rlabel metal1 3068 90 3068 100 7 nResetOut
rlabel metal1 3068 113 3068 123 7 TestOut
rlabel metal1 3068 136 3068 146 7 ClockOut
rlabel metal1 3068 159 3068 184 7 GND!
rlabel metal2 2910 0 2922 0 1 nnSDO
rlabel metal1 3068 865 3068 875 7 nSDO
rlabel metal2 216 945 228 945 5 SDO
<< end >>
