magic
tech c035u
timestamp 1384881176
<< nwell >>
rect 0 395 270 730
<< polysilicon >>
rect 44 675 51 683
rect 71 675 78 683
rect 101 675 108 683
rect 131 675 138 683
rect 44 599 51 627
rect 71 599 78 627
rect 101 599 108 627
rect 44 521 51 551
rect 71 521 78 551
rect 44 443 51 473
rect 71 443 78 473
rect 101 443 108 551
rect 44 355 51 395
rect 71 355 78 395
rect 44 295 51 325
rect 71 295 78 325
rect 101 295 108 395
rect 131 378 138 627
rect 184 482 191 490
rect 236 482 243 490
rect 184 374 191 434
rect 236 424 243 434
rect 236 410 246 424
rect 236 400 243 410
rect 239 384 243 400
rect 236 374 243 384
rect 44 215 51 265
rect 71 215 78 265
rect 101 215 108 265
rect 44 155 51 185
rect 71 155 78 185
rect 101 155 108 185
rect 131 155 138 362
rect 184 334 191 344
rect 236 336 243 344
rect 188 318 191 334
rect 44 101 51 125
rect 71 101 78 125
rect 101 101 108 125
rect 131 117 138 125
<< ndiffusion >>
rect 42 325 44 355
rect 51 325 71 355
rect 78 325 80 355
rect 41 265 44 295
rect 51 265 71 295
rect 78 265 80 295
rect 96 265 101 295
rect 108 265 110 295
rect 42 185 44 215
rect 51 185 53 215
rect 69 185 71 215
rect 78 185 80 215
rect 96 185 101 215
rect 108 185 110 215
rect 182 344 184 374
rect 191 344 218 374
rect 234 344 236 374
rect 243 344 245 374
rect 42 125 44 155
rect 51 125 71 155
rect 78 125 101 155
rect 108 125 113 155
rect 129 125 131 155
rect 138 125 140 155
<< pdiffusion >>
rect 42 627 44 675
rect 51 627 71 675
rect 78 627 80 675
rect 96 627 101 675
rect 108 627 110 675
rect 126 627 131 675
rect 138 627 140 675
rect 42 551 44 599
rect 51 551 53 599
rect 69 551 71 599
rect 78 551 80 599
rect 96 551 101 599
rect 108 551 110 599
rect 42 473 44 521
rect 51 473 53 521
rect 69 473 71 521
rect 78 473 80 521
rect 42 395 44 443
rect 51 395 71 443
rect 78 395 80 443
rect 96 395 101 443
rect 108 395 110 443
rect 182 434 184 482
rect 191 434 218 482
rect 234 434 236 482
rect 243 434 245 482
<< pohmic >>
rect 0 65 6 75
rect 22 65 34 75
rect 50 65 62 75
rect 78 65 90 75
rect 106 65 118 75
rect 134 65 146 75
rect 162 65 174 75
rect 190 65 202 75
rect 218 65 230 75
rect 246 65 270 75
<< nohmic >>
rect 0 720 6 730
rect 22 720 34 730
rect 50 720 62 730
rect 78 720 90 730
rect 106 720 118 730
rect 134 720 146 730
rect 162 720 174 730
rect 190 720 202 730
rect 218 720 230 730
rect 246 720 270 730
<< ntransistor >>
rect 44 325 51 355
rect 71 325 78 355
rect 44 265 51 295
rect 71 265 78 295
rect 101 265 108 295
rect 44 185 51 215
rect 71 185 78 215
rect 101 185 108 215
rect 184 344 191 374
rect 236 344 243 374
rect 44 125 51 155
rect 71 125 78 155
rect 101 125 108 155
rect 131 125 138 155
<< ptransistor >>
rect 44 627 51 675
rect 71 627 78 675
rect 101 627 108 675
rect 131 627 138 675
rect 44 551 51 599
rect 71 551 78 599
rect 101 551 108 599
rect 44 473 51 521
rect 71 473 78 521
rect 44 395 51 443
rect 71 395 78 443
rect 101 395 108 443
rect 184 434 191 482
rect 236 434 243 482
<< polycontact >>
rect 127 362 143 378
rect 223 384 239 400
rect 172 318 188 334
<< ndiffcontact >>
rect 26 325 42 355
rect 80 325 96 355
rect 25 265 41 295
rect 80 265 96 295
rect 110 265 126 295
rect 26 185 42 215
rect 53 185 69 215
rect 80 185 96 215
rect 110 185 126 215
rect 166 344 182 374
rect 218 344 234 374
rect 245 344 261 374
rect 26 125 42 155
rect 113 125 129 155
rect 140 125 156 155
<< pdiffcontact >>
rect 26 627 42 675
rect 80 627 96 675
rect 110 627 126 675
rect 140 627 156 675
rect 26 551 42 599
rect 53 551 69 599
rect 80 551 96 599
rect 110 551 126 599
rect 26 473 42 521
rect 53 473 69 521
rect 80 473 96 521
rect 26 395 42 443
rect 80 395 96 443
rect 110 395 126 443
rect 166 434 182 482
rect 218 434 234 482
rect 245 434 261 482
<< psubstratetap >>
rect 6 65 22 81
rect 34 65 50 81
rect 62 65 78 81
rect 90 65 106 81
rect 118 65 134 81
rect 146 65 162 81
rect 174 65 190 81
rect 202 65 218 81
rect 230 65 246 81
<< nsubstratetap >>
rect 6 714 22 730
rect 34 714 50 730
rect 62 714 78 730
rect 90 714 106 730
rect 118 714 134 730
rect 146 714 162 730
rect 174 714 190 730
rect 202 714 218 730
rect 230 714 246 730
<< metal1 >>
rect 0 760 270 770
rect 0 740 270 750
rect 0 714 6 730
rect 22 714 34 730
rect 50 714 62 730
rect 78 714 90 730
rect 106 714 118 730
rect 134 714 146 730
rect 162 714 174 730
rect 190 714 202 730
rect 218 714 230 730
rect 246 714 270 730
rect 0 705 270 714
rect 6 541 16 705
rect 29 685 208 695
rect 29 675 39 685
rect 83 675 93 685
rect 113 675 123 685
rect 29 599 39 627
rect 83 599 93 627
rect 143 580 153 627
rect 126 570 153 580
rect 56 541 66 551
rect 113 541 123 551
rect 6 531 123 541
rect 56 521 66 531
rect 96 492 116 502
rect 29 463 39 473
rect 106 463 116 492
rect 29 453 123 463
rect 29 443 39 453
rect 113 443 123 453
rect 169 403 179 434
rect 83 375 93 395
rect 198 398 208 685
rect 221 482 231 705
rect 249 424 259 434
rect 257 410 259 424
rect 29 365 127 375
rect 29 355 39 365
rect 169 374 179 389
rect 198 386 223 398
rect 143 362 146 372
rect 96 335 123 345
rect 29 315 39 325
rect 29 305 93 315
rect 29 295 39 305
rect 83 295 93 305
rect 113 295 123 335
rect 136 330 146 362
rect 136 320 172 330
rect 113 255 123 265
rect 6 245 123 255
rect 6 90 16 245
rect 198 235 208 386
rect 249 374 259 410
rect 29 225 208 235
rect 29 215 39 225
rect 83 215 93 225
rect 29 155 39 185
rect 56 175 66 185
rect 113 175 123 185
rect 56 165 153 175
rect 143 155 153 165
rect 119 90 129 125
rect 221 90 231 344
rect 0 81 270 90
rect 0 65 6 81
rect 22 65 34 81
rect 50 65 62 81
rect 78 65 90 81
rect 106 65 118 81
rect 134 65 146 81
rect 162 65 174 81
rect 190 65 202 81
rect 218 65 230 81
rect 246 65 270 81
rect 0 45 270 55
rect 0 25 270 35
rect 0 5 270 15
<< m2contact >>
rect 166 389 180 403
rect 243 410 257 424
rect 44 101 58 115
rect 70 101 84 115
rect 94 101 108 115
<< metal2 >>
rect 48 115 60 775
rect 72 115 84 775
rect 96 115 108 775
rect 168 403 180 775
rect 58 101 60 115
rect 48 0 60 101
rect 72 0 84 101
rect 96 0 108 101
rect 168 0 180 389
rect 240 424 252 775
rect 240 410 243 424
rect 240 0 252 410
<< labels >>
rlabel metal1 0 65 0 90 3 GND!
rlabel metal1 270 65 270 90 7 GND!
rlabel metal1 270 705 270 730 7 Vdd!
rlabel metal1 0 705 0 730 3 Vdd!
rlabel metal1 0 740 0 750 3 Q
rlabel metal1 0 760 0 770 3 ScanReturn
rlabel metal1 270 760 270 770 7 ScanReturn
rlabel metal1 270 740 270 750 7 Q
rlabel metal1 0 25 0 35 3 Test
rlabel metal1 0 45 0 55 3 Clock
rlabel metal1 270 25 270 35 7 Test
rlabel metal1 270 45 270 55 7 Clock
rlabel metal2 48 0 60 0 1 A
rlabel metal2 72 0 84 0 1 B
rlabel metal2 96 0 108 0 1 Cin
rlabel metal2 168 0 180 0 1 Cout
rlabel metal2 240 0 252 0 1 S
rlabel metal1 0 5 0 15 3 Reset
rlabel metal1 270 5 270 15 7 Reset
rlabel metal2 48 775 60 775 5 A
rlabel metal2 72 775 84 775 5 B
rlabel metal2 96 775 108 775 5 Cin
rlabel metal2 168 775 180 775 5 Cout
rlabel metal2 240 775 252 775 5 S
<< end >>
