magic
tech c035u
timestamp 1386275188
<< metal1 >>
rect 6 833 250 843
rect 6 769 16 833
rect 43 792 53 809
rect 32 782 59 792
rect 0 759 59 769
rect 0 721 59 746
<< m2contact >>
rect 250 831 264 845
rect 41 809 55 823
<< metal2 >>
rect 83 821 95 858
rect 55 809 95 821
rect 83 799 95 809
rect 203 799 215 858
rect 251 799 263 831
use inv inv_1
timestamp 1386238110
transform 1 0 59 0 1 0
box 0 0 120 799
use inv inv_0
timestamp 1386238110
transform 1 0 179 0 1 0
box 0 0 120 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 299 0 1 0
box 0 0 320 799
<< labels >>
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 759 0 769 3 Scan
rlabel metal2 203 858 215 858 5 ScanIn
rlabel metal2 83 858 95 858 5 nScan
<< end >>
