magic
tech c035u
timestamp 1385906230
<< nwell >>
rect 0 302 360 646
<< polysilicon >>
rect 44 572 49 585
rect 73 572 78 585
rect 44 531 51 572
rect 71 531 78 572
rect 91 531 98 595
rect 118 531 125 572
rect 148 531 155 570
rect 175 531 182 572
rect 206 531 213 595
rect 279 531 286 539
rect 44 404 51 483
rect 71 404 78 483
rect 91 404 98 483
rect 118 404 125 483
rect 44 261 51 356
rect 71 261 78 356
rect 91 261 98 356
rect 118 261 125 356
rect 148 287 155 483
rect 44 161 51 231
rect 71 161 78 231
rect 91 161 98 231
rect 118 161 125 231
rect 148 161 155 271
rect 175 161 182 483
rect 206 404 213 483
rect 279 450 286 484
rect 269 443 286 450
rect 206 261 213 356
rect 206 161 213 231
rect 262 207 269 437
rect 292 404 299 412
rect 292 287 299 356
rect 292 261 299 271
rect 292 223 299 231
rect 262 161 269 191
rect 44 123 51 131
rect 71 123 78 131
rect 91 123 98 131
rect 118 123 125 131
rect 148 123 155 131
rect 175 123 182 131
rect 206 123 213 131
rect 262 123 269 131
<< ndiffusion >>
rect 42 231 44 261
rect 51 231 53 261
rect 69 231 71 261
rect 78 231 91 261
rect 98 231 100 261
rect 116 231 118 261
rect 125 231 127 261
rect 204 231 206 261
rect 213 231 215 261
rect 290 231 292 261
rect 299 231 301 261
rect 42 131 44 161
rect 51 131 53 161
rect 69 131 71 161
rect 78 131 91 161
rect 98 131 118 161
rect 125 131 127 161
rect 143 131 148 161
rect 155 131 157 161
rect 173 131 175 161
rect 182 131 188 161
rect 204 131 206 161
rect 213 131 215 161
rect 260 131 262 161
rect 269 131 271 161
<< pdiffusion >>
rect 42 483 44 531
rect 51 483 53 531
rect 69 483 71 531
rect 78 483 91 531
rect 98 483 118 531
rect 125 483 127 531
rect 143 483 148 531
rect 155 483 157 531
rect 173 483 175 531
rect 182 483 188 531
rect 204 483 206 531
rect 213 483 215 531
rect 277 484 279 531
rect 286 484 288 531
rect 42 356 44 404
rect 51 356 53 404
rect 69 356 71 404
rect 78 356 91 404
rect 98 356 100 404
rect 116 356 118 404
rect 125 356 127 404
rect 204 356 206 404
rect 213 356 215 404
rect 290 356 292 404
rect 299 356 301 404
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 174 86
rect 190 76 202 86
rect 218 76 230 86
rect 246 76 258 86
rect 274 76 286 86
rect 302 76 314 86
rect 330 76 360 86
<< nohmic >>
rect 0 636 6 646
rect 22 636 34 646
rect 50 636 62 646
rect 78 636 90 646
rect 106 636 118 646
rect 134 636 146 646
rect 162 636 174 646
rect 190 636 202 646
rect 218 636 230 646
rect 246 636 258 646
rect 274 636 286 646
rect 302 636 314 646
rect 330 636 360 646
<< ntransistor >>
rect 44 231 51 261
rect 71 231 78 261
rect 91 231 98 261
rect 118 231 125 261
rect 206 231 213 261
rect 292 231 299 261
rect 44 131 51 161
rect 71 131 78 161
rect 91 131 98 161
rect 118 131 125 161
rect 148 131 155 161
rect 175 131 182 161
rect 206 131 213 161
rect 262 131 269 161
<< ptransistor >>
rect 44 483 51 531
rect 71 483 78 531
rect 91 483 98 531
rect 118 483 125 531
rect 148 483 155 531
rect 175 483 182 531
rect 206 483 213 531
rect 279 484 286 531
rect 44 356 51 404
rect 71 356 78 404
rect 91 356 98 404
rect 118 356 125 404
rect 206 356 213 404
rect 292 356 299 404
<< polycontact >>
rect 87 595 103 611
rect 202 595 218 611
rect 49 572 73 588
rect 113 572 129 588
rect 166 572 182 588
rect 143 271 159 287
rect 253 437 269 453
rect 288 271 304 287
rect 253 191 269 207
<< ndiffcontact >>
rect 26 231 42 261
rect 53 231 69 261
rect 100 231 116 261
rect 127 231 143 261
rect 188 231 204 261
rect 215 231 231 261
rect 274 231 290 261
rect 301 231 317 261
rect 26 131 42 161
rect 53 131 69 161
rect 127 131 143 161
rect 157 131 173 161
rect 188 131 204 161
rect 215 131 231 161
rect 244 131 260 161
rect 271 131 287 161
<< pdiffcontact >>
rect 26 483 42 531
rect 53 483 69 531
rect 127 483 143 531
rect 157 483 173 531
rect 188 483 204 531
rect 215 483 231 531
rect 261 484 277 531
rect 288 484 304 531
rect 26 356 42 404
rect 53 356 69 404
rect 100 356 116 404
rect 127 356 143 404
rect 188 356 204 404
rect 215 356 231 404
rect 274 356 290 404
rect 301 356 317 404
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
rect 174 76 190 92
rect 202 76 218 92
rect 230 76 246 92
rect 258 76 274 92
rect 286 76 302 92
rect 314 76 330 92
<< nsubstratetap >>
rect 6 630 22 646
rect 34 630 50 646
rect 62 630 78 646
rect 90 630 106 646
rect 118 630 134 646
rect 146 630 162 646
rect 174 630 190 646
rect 202 630 218 646
rect 230 630 246 646
rect 258 630 274 646
rect 286 630 302 646
rect 314 630 330 646
<< metal1 >>
rect 0 682 360 692
rect 0 659 360 669
rect 0 630 6 646
rect 22 630 34 646
rect 50 630 62 646
rect 78 630 90 646
rect 106 630 118 646
rect 134 630 146 646
rect 162 630 174 646
rect 190 630 202 646
rect 218 630 230 646
rect 246 630 258 646
rect 274 630 286 646
rect 302 630 314 646
rect 330 630 360 646
rect 0 621 360 630
rect 29 531 39 621
rect 49 588 63 597
rect 103 598 139 608
rect 153 598 202 608
rect 129 575 142 585
rect 156 575 166 585
rect 56 541 228 551
rect 56 531 66 541
rect 160 531 170 541
rect 218 531 228 541
rect 29 404 39 483
rect 129 453 141 483
rect 191 473 201 483
rect 241 473 251 621
rect 264 531 274 569
rect 294 531 304 621
rect 191 463 251 473
rect 129 441 253 453
rect 291 424 301 484
rect 56 414 140 424
rect 56 404 66 414
rect 130 404 140 414
rect 280 414 301 424
rect 280 404 290 414
rect 143 375 188 385
rect 231 374 274 384
rect 103 281 113 356
rect 317 288 327 366
rect 6 271 66 281
rect 6 101 16 271
rect 56 261 66 271
rect 103 271 143 281
rect 159 271 288 281
rect 103 261 113 271
rect 143 242 188 252
rect 231 241 274 251
rect 317 251 327 274
rect 29 221 39 231
rect 130 221 140 231
rect 29 211 140 221
rect 56 191 253 201
rect 56 161 66 191
rect 107 171 170 181
rect 29 121 39 131
rect 107 121 117 171
rect 160 161 170 171
rect 191 161 201 191
rect 279 181 289 231
rect 277 171 289 181
rect 244 161 257 167
rect 277 161 287 171
rect 29 111 117 121
rect 130 101 140 131
rect 160 121 170 131
rect 218 121 228 131
rect 160 111 228 121
rect 274 101 284 131
rect 0 92 360 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 174 92
rect 190 76 202 92
rect 218 76 230 92
rect 246 76 258 92
rect 274 76 286 92
rect 302 76 314 92
rect 330 76 360 92
rect 0 53 360 63
rect 0 30 360 40
rect 0 7 360 17
<< m2contact >>
rect 49 597 63 611
rect 139 597 153 611
rect 142 573 156 587
rect 262 569 276 583
rect 316 274 330 288
rect 241 167 255 181
<< metal2 >>
rect 48 611 60 699
rect 120 611 132 699
rect 48 597 49 611
rect 120 597 139 611
rect 48 0 60 597
rect 120 0 132 597
rect 168 587 180 699
rect 156 573 180 587
rect 168 0 180 573
rect 240 582 252 699
rect 240 570 262 582
rect 240 181 252 570
rect 312 288 324 699
rect 312 274 316 288
rect 240 167 241 181
rect 240 0 252 167
rect 312 0 324 274
<< labels >>
rlabel metal1 360 53 360 63 7 Clock
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 360 76 360 101 7 GND!
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 360 30 360 40 7 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal2 48 0 60 0 1 A
rlabel metal2 120 0 132 0 1 B
rlabel metal2 168 0 180 0 1 Cin
rlabel metal2 312 0 324 0 1 Cout
rlabel metal2 240 0 252 0 1 S
rlabel metal1 360 7 360 17 8 nReset
rlabel metal1 0 659 0 669 3 Scan
rlabel metal1 360 659 360 669 7 Scan
rlabel metal2 168 699 180 699 5 Cin
rlabel metal2 120 699 132 699 5 B
rlabel metal2 48 699 60 699 5 A
rlabel metal1 0 682 0 692 3 ScanReturn
rlabel metal2 240 699 252 699 5 S
rlabel metal2 312 699 324 699 5 Cout
rlabel metal1 360 682 360 692 7 ScanReturn
rlabel metal1 0 621 0 646 3 Vdd!
rlabel metal1 360 621 360 646 7 Vdd!
<< end >>
