magic
tech c035u
timestamp 1385926557
<< nwell >>
rect 202 392 1464 736
rect 405 391 451 392
rect 742 391 788 392
rect 1079 391 1125 392
<< polysilicon >>
rect 538 682 545 690
rect 565 682 572 690
rect 592 682 599 690
rect 619 682 626 690
rect 875 682 882 690
rect 902 682 909 690
rect 929 682 936 690
rect 956 682 963 690
rect 1212 682 1219 690
rect 1239 682 1246 690
rect 1266 682 1273 690
rect 1293 682 1300 690
rect 480 604 487 612
rect 507 604 514 612
rect 425 549 432 557
rect 370 450 377 458
rect 817 604 824 612
rect 844 604 851 612
rect 762 549 769 557
rect 707 450 714 458
rect 1154 604 1161 612
rect 1181 604 1188 612
rect 1099 549 1106 557
rect 1044 450 1051 458
rect 1394 506 1396 522
rect 1389 461 1396 506
rect 370 378 377 392
rect 425 378 432 392
rect 480 379 487 392
rect 375 362 377 378
rect 430 362 432 378
rect 485 375 487 379
rect 507 375 514 392
rect 538 379 545 392
rect 485 368 514 375
rect 485 363 487 368
rect 543 375 545 379
rect 565 375 572 392
rect 592 375 599 392
rect 619 375 626 392
rect 707 378 714 392
rect 762 378 769 392
rect 817 379 824 392
rect 543 368 626 375
rect 543 363 545 368
rect 370 352 377 362
rect 425 352 432 362
rect 480 352 487 363
rect 538 352 545 363
rect 565 352 572 368
rect 712 362 714 378
rect 767 362 769 378
rect 822 375 824 379
rect 844 375 851 392
rect 875 379 882 392
rect 822 368 851 375
rect 822 363 824 368
rect 880 375 882 379
rect 902 375 909 392
rect 929 375 936 392
rect 956 375 963 392
rect 1044 378 1051 392
rect 1099 378 1106 392
rect 1154 379 1161 392
rect 880 368 963 375
rect 880 363 882 368
rect 707 352 714 362
rect 762 352 769 362
rect 817 352 824 363
rect 875 352 882 363
rect 902 352 909 368
rect 1049 362 1051 378
rect 1104 362 1106 378
rect 1159 375 1161 379
rect 1181 375 1188 392
rect 1212 379 1219 392
rect 1159 368 1188 375
rect 1159 363 1161 368
rect 1217 375 1219 379
rect 1239 375 1246 392
rect 1266 375 1273 392
rect 1293 375 1300 392
rect 1217 368 1300 375
rect 1217 363 1219 368
rect 1044 352 1051 362
rect 1099 352 1106 362
rect 1154 352 1161 363
rect 1212 352 1219 363
rect 1239 352 1246 368
rect 1389 367 1396 413
rect 370 324 377 332
rect 425 290 432 298
rect 480 198 487 206
rect 707 324 714 332
rect 762 290 769 298
rect 817 198 824 206
rect 1044 324 1051 332
rect 1099 290 1106 298
rect 1154 198 1161 206
rect 1389 329 1396 337
rect 538 144 545 152
rect 565 144 572 152
rect 875 144 882 152
rect 902 144 909 152
rect 1212 144 1219 152
rect 1239 144 1246 152
<< ndiffusion >>
rect 368 332 370 352
rect 377 332 379 352
rect 423 298 425 352
rect 432 298 434 352
rect 478 206 480 352
rect 487 206 489 352
rect 536 152 538 352
rect 545 152 547 352
rect 563 152 565 352
rect 572 152 574 352
rect 705 332 707 352
rect 714 332 716 352
rect 760 298 762 352
rect 769 298 771 352
rect 815 206 817 352
rect 824 206 826 352
rect 873 152 875 352
rect 882 152 884 352
rect 900 152 902 352
rect 909 152 911 352
rect 1042 332 1044 352
rect 1051 332 1053 352
rect 1097 298 1099 352
rect 1106 298 1108 352
rect 1152 206 1154 352
rect 1161 206 1163 352
rect 1210 152 1212 352
rect 1219 152 1221 352
rect 1237 152 1239 352
rect 1246 152 1248 352
rect 1387 337 1389 367
rect 1396 337 1398 367
<< pdiffusion >>
rect 368 392 370 450
rect 377 392 379 450
rect 423 392 425 549
rect 432 392 434 549
rect 478 392 480 604
rect 487 392 489 604
rect 505 392 507 604
rect 514 392 516 604
rect 536 392 538 682
rect 545 392 547 682
rect 563 392 565 682
rect 572 392 574 682
rect 590 392 592 682
rect 599 392 601 682
rect 617 392 619 682
rect 626 392 628 682
rect 705 392 707 450
rect 714 392 716 450
rect 760 392 762 549
rect 769 392 771 549
rect 815 392 817 604
rect 824 392 826 604
rect 842 392 844 604
rect 851 392 853 604
rect 873 392 875 682
rect 882 392 884 682
rect 900 392 902 682
rect 909 392 911 682
rect 927 392 929 682
rect 936 392 938 682
rect 954 392 956 682
rect 963 392 965 682
rect 1042 392 1044 450
rect 1051 392 1053 450
rect 1097 392 1099 549
rect 1106 392 1108 549
rect 1152 392 1154 604
rect 1161 392 1163 604
rect 1179 392 1181 604
rect 1188 392 1190 604
rect 1210 392 1212 682
rect 1219 392 1221 682
rect 1237 392 1239 682
rect 1246 392 1248 682
rect 1264 392 1266 682
rect 1273 392 1275 682
rect 1291 392 1293 682
rect 1300 392 1302 682
rect 1387 413 1389 461
rect 1396 413 1398 461
<< pohmic >>
rect 320 66 326 76
rect 342 66 354 76
rect 370 66 382 76
rect 398 66 410 76
rect 426 66 438 76
rect 454 66 466 76
rect 482 66 494 76
rect 510 66 522 76
rect 538 66 550 76
rect 567 66 579 76
rect 595 66 607 76
rect 623 66 635 76
rect 651 66 663 76
rect 679 66 691 76
rect 707 66 719 76
rect 735 66 747 76
rect 763 66 775 76
rect 791 66 803 76
rect 819 66 831 76
rect 847 66 859 76
rect 875 66 887 76
rect 904 66 916 76
rect 932 66 944 76
rect 960 66 972 76
rect 988 66 1000 76
rect 1016 66 1028 76
rect 1044 66 1056 76
rect 1072 66 1084 76
rect 1100 66 1112 76
rect 1128 66 1140 76
rect 1156 66 1168 76
rect 1184 66 1196 76
rect 1212 66 1224 76
rect 1241 66 1253 76
rect 1269 66 1281 76
rect 1297 66 1309 76
rect 1325 66 1337 76
rect 1353 66 1365 76
rect 1381 66 1393 76
rect 1409 66 1421 76
rect 1437 66 1464 76
<< nohmic >>
rect 202 726 214 736
rect 230 726 242 736
rect 258 726 270 736
rect 286 726 298 736
rect 314 726 326 736
rect 342 726 354 736
rect 370 726 382 736
rect 398 726 410 736
rect 426 726 438 736
rect 454 726 466 736
rect 482 726 494 736
rect 510 726 522 736
rect 538 726 550 736
rect 567 726 579 736
rect 595 726 607 736
rect 623 726 635 736
rect 651 726 663 736
rect 679 726 691 736
rect 707 726 719 736
rect 735 726 747 736
rect 763 726 775 736
rect 791 726 803 736
rect 819 726 831 736
rect 847 726 859 736
rect 875 726 887 736
rect 904 726 916 736
rect 932 726 944 736
rect 960 726 972 736
rect 988 726 1000 736
rect 1016 726 1028 736
rect 1044 726 1056 736
rect 1072 726 1084 736
rect 1100 726 1112 736
rect 1128 726 1140 736
rect 1156 726 1168 736
rect 1184 726 1196 736
rect 1212 726 1224 736
rect 1241 726 1253 736
rect 1269 726 1281 736
rect 1297 726 1309 736
rect 1325 726 1337 736
rect 1353 726 1365 736
rect 1381 726 1393 736
rect 1409 726 1421 736
rect 1437 726 1464 736
<< ntransistor >>
rect 370 332 377 352
rect 425 298 432 352
rect 480 206 487 352
rect 538 152 545 352
rect 565 152 572 352
rect 707 332 714 352
rect 762 298 769 352
rect 817 206 824 352
rect 875 152 882 352
rect 902 152 909 352
rect 1044 332 1051 352
rect 1099 298 1106 352
rect 1154 206 1161 352
rect 1212 152 1219 352
rect 1239 152 1246 352
rect 1389 337 1396 367
<< ptransistor >>
rect 370 392 377 450
rect 425 392 432 549
rect 480 392 487 604
rect 507 392 514 604
rect 538 392 545 682
rect 565 392 572 682
rect 592 392 599 682
rect 619 392 626 682
rect 707 392 714 450
rect 762 392 769 549
rect 817 392 824 604
rect 844 392 851 604
rect 875 392 882 682
rect 902 392 909 682
rect 929 392 936 682
rect 956 392 963 682
rect 1044 392 1051 450
rect 1099 392 1106 549
rect 1154 392 1161 604
rect 1181 392 1188 604
rect 1212 392 1219 682
rect 1239 392 1246 682
rect 1266 392 1273 682
rect 1293 392 1300 682
rect 1389 413 1396 461
<< polycontact >>
rect 1378 506 1394 522
rect 359 362 375 378
rect 414 362 430 378
rect 469 363 485 379
rect 527 363 543 379
rect 696 362 712 378
rect 751 362 767 378
rect 806 363 822 379
rect 864 363 880 379
rect 1033 362 1049 378
rect 1088 362 1104 378
rect 1143 363 1159 379
rect 1201 363 1217 379
<< ndiffcontact >>
rect 352 332 368 352
rect 379 332 395 352
rect 407 298 423 352
rect 434 298 450 352
rect 462 206 478 352
rect 489 206 505 352
rect 520 152 536 352
rect 547 152 563 352
rect 574 152 590 352
rect 689 332 705 352
rect 716 332 732 352
rect 744 298 760 352
rect 771 298 787 352
rect 799 206 815 352
rect 826 206 842 352
rect 857 152 873 352
rect 884 152 900 352
rect 911 152 927 352
rect 1026 332 1042 352
rect 1053 332 1069 352
rect 1081 298 1097 352
rect 1108 298 1124 352
rect 1136 206 1152 352
rect 1163 206 1179 352
rect 1194 152 1210 352
rect 1221 152 1237 352
rect 1248 152 1264 352
rect 1371 337 1387 367
rect 1398 337 1414 367
<< pdiffcontact >>
rect 519 604 536 682
rect 352 392 368 450
rect 379 392 395 450
rect 407 392 423 549
rect 434 392 450 549
rect 462 392 478 604
rect 489 392 505 604
rect 516 392 536 604
rect 547 392 563 682
rect 574 392 590 682
rect 601 392 617 682
rect 628 392 644 682
rect 856 604 873 682
rect 689 392 705 450
rect 716 392 732 450
rect 744 392 760 549
rect 771 392 787 549
rect 799 392 815 604
rect 826 392 842 604
rect 853 392 873 604
rect 884 392 900 682
rect 911 392 927 682
rect 938 392 954 682
rect 965 392 981 682
rect 1193 604 1210 682
rect 1026 392 1042 450
rect 1053 392 1069 450
rect 1081 392 1097 549
rect 1108 392 1124 549
rect 1136 392 1152 604
rect 1163 392 1179 604
rect 1190 392 1210 604
rect 1221 392 1237 682
rect 1248 392 1264 682
rect 1275 392 1291 682
rect 1302 392 1318 682
rect 1371 413 1387 461
rect 1398 413 1414 461
<< psubstratetap >>
rect 326 66 342 82
rect 354 66 370 82
rect 382 66 398 82
rect 410 66 426 82
rect 438 66 454 82
rect 466 66 482 82
rect 494 66 510 82
rect 522 66 538 82
rect 550 66 567 82
rect 579 66 595 82
rect 607 66 623 82
rect 635 66 651 82
rect 663 66 679 82
rect 691 66 707 82
rect 719 66 735 82
rect 747 66 763 82
rect 775 66 791 82
rect 803 66 819 82
rect 831 66 847 82
rect 859 66 875 82
rect 887 66 904 82
rect 916 66 932 82
rect 944 66 960 82
rect 972 66 988 82
rect 1000 66 1016 82
rect 1028 66 1044 82
rect 1056 66 1072 82
rect 1084 66 1100 82
rect 1112 66 1128 82
rect 1140 66 1156 82
rect 1168 66 1184 82
rect 1196 66 1212 82
rect 1224 66 1241 82
rect 1253 66 1269 82
rect 1281 66 1297 82
rect 1309 66 1325 82
rect 1337 66 1353 82
rect 1365 66 1381 82
rect 1393 66 1409 82
rect 1421 66 1437 82
<< nsubstratetap >>
rect 214 720 230 736
rect 242 720 258 736
rect 270 720 286 736
rect 298 720 314 736
rect 326 720 342 736
rect 354 720 370 736
rect 382 720 398 736
rect 410 720 426 736
rect 438 720 454 736
rect 466 720 482 736
rect 494 720 510 736
rect 522 720 538 736
rect 550 720 567 736
rect 579 720 595 736
rect 607 720 623 736
rect 635 720 651 736
rect 663 720 679 736
rect 691 720 707 736
rect 719 720 735 736
rect 747 720 763 736
rect 775 720 791 736
rect 803 720 819 736
rect 831 720 847 736
rect 859 720 875 736
rect 887 720 904 736
rect 916 720 932 736
rect 944 720 960 736
rect 972 720 988 736
rect 1000 720 1016 736
rect 1028 720 1044 736
rect 1056 720 1072 736
rect 1084 720 1100 736
rect 1112 720 1128 736
rect 1140 720 1156 736
rect 1168 720 1184 736
rect 1196 720 1212 736
rect 1224 720 1241 736
rect 1253 720 1269 736
rect 1281 720 1297 736
rect 1309 720 1325 736
rect 1337 720 1353 736
rect 1365 720 1381 736
rect 1393 720 1409 736
rect 1421 720 1437 736
<< metal1 >>
rect 190 749 200 782
rect 229 772 1356 782
rect 1400 772 1464 782
rect 229 749 1464 759
rect 200 720 214 736
rect 230 720 242 736
rect 258 720 270 736
rect 286 720 298 736
rect 314 720 326 736
rect 342 720 354 736
rect 370 720 382 736
rect 398 720 410 736
rect 426 720 438 736
rect 454 720 466 736
rect 482 720 494 736
rect 510 720 522 736
rect 538 720 550 736
rect 567 720 579 736
rect 595 720 607 736
rect 623 720 635 736
rect 651 720 663 736
rect 679 720 691 736
rect 707 720 719 736
rect 735 720 747 736
rect 763 720 775 736
rect 791 720 803 736
rect 819 720 831 736
rect 847 720 859 736
rect 875 720 887 736
rect 904 720 916 736
rect 932 720 944 736
rect 960 720 972 736
rect 988 720 1000 736
rect 1016 720 1028 736
rect 1044 720 1056 736
rect 1072 720 1084 736
rect 1100 720 1112 736
rect 1128 720 1140 736
rect 1156 720 1168 736
rect 1184 720 1196 736
rect 1212 720 1224 736
rect 1241 720 1253 736
rect 1269 720 1281 736
rect 1297 720 1309 736
rect 1325 720 1337 736
rect 1353 720 1365 736
rect 1381 720 1393 736
rect 1409 720 1421 736
rect 1437 720 1464 736
rect 200 711 1464 720
rect 352 450 368 711
rect 407 549 423 711
rect 462 604 478 711
rect 516 682 536 711
rect 574 682 590 711
rect 628 682 644 711
rect 516 604 519 682
rect 689 450 705 711
rect 744 549 760 711
rect 799 604 815 711
rect 853 682 873 711
rect 911 682 927 711
rect 965 682 981 711
rect 853 604 856 682
rect 1026 450 1042 711
rect 1081 549 1097 711
rect 1136 604 1152 711
rect 1190 682 1210 711
rect 1248 682 1264 711
rect 1302 682 1318 711
rect 1190 604 1193 682
rect 1380 522 1394 528
rect 1404 461 1414 711
rect 240 340 252 377
rect 277 365 359 375
rect 263 353 277 363
rect 385 375 395 392
rect 385 365 414 375
rect 385 352 395 365
rect 440 376 450 392
rect 440 366 469 376
rect 440 352 450 366
rect 495 376 505 392
rect 495 366 527 376
rect 495 352 505 366
rect 553 377 563 392
rect 607 379 617 392
rect 553 367 606 377
rect 553 352 563 367
rect 667 365 696 375
rect 722 375 732 392
rect 722 365 751 375
rect 722 352 732 365
rect 777 376 787 392
rect 777 366 806 376
rect 777 352 787 366
rect 832 376 842 392
rect 832 366 864 376
rect 832 352 842 366
rect 890 377 900 392
rect 944 379 954 392
rect 890 367 944 377
rect 890 352 900 367
rect 1022 365 1033 375
rect 1059 375 1069 392
rect 1059 365 1088 375
rect 1059 352 1069 365
rect 1114 376 1124 392
rect 1114 366 1143 376
rect 1114 352 1124 366
rect 1169 376 1179 392
rect 1169 366 1201 376
rect 1169 352 1179 366
rect 1227 377 1237 392
rect 1281 379 1291 392
rect 1227 367 1279 377
rect 1227 352 1237 367
rect 1371 367 1381 413
rect 352 91 368 332
rect 407 91 423 298
rect 462 91 478 206
rect 520 91 536 152
rect 574 91 590 152
rect 689 91 705 332
rect 744 91 760 298
rect 799 91 815 206
rect 857 91 873 152
rect 911 91 927 152
rect 1026 91 1042 332
rect 1081 91 1097 298
rect 1136 91 1152 206
rect 1194 91 1210 152
rect 1248 91 1264 152
rect 1398 91 1408 337
rect 320 82 1464 91
rect 320 66 326 82
rect 342 66 354 82
rect 370 66 382 82
rect 398 66 410 82
rect 426 66 438 82
rect 454 66 466 82
rect 482 66 494 82
rect 510 66 522 82
rect 538 66 550 82
rect 567 66 579 82
rect 595 66 607 82
rect 623 66 635 82
rect 651 66 663 82
rect 679 66 691 82
rect 707 66 719 82
rect 735 66 747 82
rect 763 66 775 82
rect 791 66 803 82
rect 819 66 831 82
rect 847 66 859 82
rect 875 66 887 82
rect 904 66 916 82
rect 932 66 944 82
rect 960 66 972 82
rect 988 66 1000 82
rect 1016 66 1028 82
rect 1044 66 1056 82
rect 1072 66 1084 82
rect 1100 66 1112 82
rect 1128 66 1140 82
rect 1156 66 1168 82
rect 1184 66 1196 82
rect 1212 66 1224 82
rect 1241 66 1253 82
rect 1269 66 1281 82
rect 1297 66 1309 82
rect 1325 66 1337 82
rect 1353 66 1365 82
rect 1381 66 1393 82
rect 1409 66 1421 82
rect 1437 66 1464 82
rect 216 -3 228 56
rect 239 33 253 43
rect 620 43 1464 53
rect 253 20 653 30
rect 959 20 1464 30
rect 301 -3 1009 7
rect 1033 -3 1270 7
rect 1294 -3 1304 7
rect 1318 -3 1464 7
<< m2contact >>
rect 215 770 229 784
rect 1356 771 1370 785
rect 1386 771 1400 785
rect 215 746 229 760
rect 0 711 200 736
rect 1380 528 1394 542
rect 1357 447 1371 461
rect 263 363 277 377
rect 263 339 277 353
rect 606 365 620 379
rect 653 363 667 377
rect 944 365 958 379
rect 1008 363 1022 377
rect 1279 365 1293 379
rect 239 43 253 57
rect 606 41 620 55
rect 239 19 253 33
rect 653 18 667 32
rect 945 19 959 33
rect 239 -5 253 9
rect 263 -5 277 9
rect 287 -5 301 9
rect 1009 -5 1023 9
rect 1280 -5 1294 9
rect 1304 -5 1318 9
<< metal2 >>
rect 0 736 200 789
rect 216 784 228 789
rect 0 -10 200 711
rect 216 -10 228 746
rect 240 57 252 789
rect 264 377 276 789
rect 264 353 276 363
rect 240 33 252 43
rect 240 9 252 19
rect 264 9 276 339
rect 288 9 300 789
rect 1358 461 1370 771
rect 1386 542 1398 771
rect 1394 528 1398 542
rect 607 55 619 365
rect 654 32 666 363
rect 946 33 958 365
rect 1010 9 1022 363
rect 1281 9 1293 365
rect 1294 -5 1304 9
rect 240 -10 252 -5
rect 264 -10 276 -5
rect 288 -10 300 -5
<< labels >>
rlabel metal2 0 789 200 789 5 Vdd!
rlabel metal2 0 -10 200 -10 1 Vdd!
rlabel metal1 1464 711 1464 736 7 Vdd!
rlabel metal1 1464 749 1464 759 7 SDI
rlabel metal1 1464 772 1464 782 7 nSDO
rlabel metal1 1464 43 1464 53 7 ClockOut
rlabel metal1 1464 20 1464 30 7 TestOut
rlabel metal1 1464 -3 1464 7 7 nResetOut
rlabel metal1 1464 66 1464 91 7 GND!
rlabel metal2 216 -10 228 -10 1 SDI
rlabel metal2 240 -10 252 -10 1 Test
rlabel metal2 264 -10 276 -10 1 Clock
rlabel metal2 288 -10 300 -10 1 nReset
rlabel metal2 288 789 300 789 5 nReset
rlabel metal2 240 789 252 789 5 Test
rlabel metal2 264 789 276 789 5 Clock
rlabel metal2 216 789 228 789 5 SDO
<< end >>
