magic
tech c035u
timestamp 1385031732
<< nwell >>
rect 0 522 116 734
<< polysilicon >>
rect 55 570 62 578
rect 55 511 62 522
rect 60 495 62 511
rect 55 482 62 495
rect 55 444 62 452
<< ndiffusion >>
rect 53 452 55 482
rect 62 452 64 482
<< pdiffusion >>
rect 53 522 55 570
rect 62 522 64 570
<< pohmic >>
rect 0 74 6 84
rect 22 74 34 84
rect 50 74 62 84
rect 78 74 90 84
rect 106 74 116 84
<< nohmic >>
rect 0 724 6 734
rect 22 724 34 734
rect 50 724 62 734
rect 78 724 90 734
rect 106 724 116 734
<< ntransistor >>
rect 55 452 62 482
<< ptransistor >>
rect 55 522 62 570
<< polycontact >>
rect 44 495 60 511
<< ndiffcontact >>
rect 37 452 53 482
rect 64 452 80 482
<< pdiffcontact >>
rect 37 522 53 570
rect 64 522 80 570
<< psubstratetap >>
rect 6 74 22 90
rect 34 74 50 90
rect 62 74 78 90
rect 90 74 106 90
<< nsubstratetap >>
rect 6 718 22 734
rect 34 718 50 734
rect 62 718 78 734
rect 90 718 106 734
<< metal1 >>
rect 0 770 116 780
rect 0 747 116 757
rect 0 718 6 734
rect 22 718 34 734
rect 50 718 62 734
rect 78 718 90 734
rect 106 718 116 734
rect 0 709 116 718
rect 37 570 53 709
rect 34 498 44 508
rect 70 509 80 522
rect 70 482 80 495
rect 36 99 52 452
rect 0 90 116 99
rect 0 74 6 90
rect 22 74 34 90
rect 50 74 62 90
rect 78 74 90 90
rect 106 74 116 90
rect 0 51 116 61
rect 0 28 116 38
rect 0 5 116 15
<< m2contact >>
rect 20 496 34 510
rect 70 495 84 509
<< metal2 >>
rect 24 510 36 785
rect 34 496 36 510
rect 72 509 84 785
rect 24 0 36 496
rect 72 0 84 495
<< labels >>
rlabel metal1 116 5 116 15 8 nReset
rlabel metal1 116 28 116 38 7 Test
rlabel metal1 116 51 116 61 7 Clock
rlabel metal1 116 74 116 99 7 GND!
rlabel metal1 116 709 116 734 7 Vdd!
rlabel metal1 116 747 116 757 7 Scan
rlabel metal1 116 770 116 780 6 ScanReturn
rlabel metal2 24 0 36 0 1 A
rlabel metal2 24 785 36 785 5 A
rlabel metal2 72 785 84 785 5 Y
rlabel metal2 72 0 84 0 1 Y
rlabel metal1 0 74 0 99 7 GND!
rlabel metal1 0 51 0 61 7 Clock
rlabel metal1 0 28 0 38 7 Test
rlabel metal1 0 5 0 15 8 nReset
rlabel metal1 0 709 0 734 7 Vdd!
rlabel metal1 0 747 0 757 7 Scan
rlabel metal1 0 770 0 780 6 ScanReturn
<< end >>
