magic
tech c035u
timestamp 1384964622
<< error_p >>
rect 23 194 24 195
<< nwell >>
rect 0 128 99 217
<< polysilicon >>
rect 28 183 35 191
rect 55 183 62 191
rect 28 3 35 135
rect 55 65 62 135
rect 61 49 62 65
rect 28 -23 35 -13
rect 55 -23 62 49
rect 28 -61 35 -53
rect 55 -61 62 -53
<< ndiffusion >>
rect 26 -53 28 -23
rect 35 -53 55 -23
rect 62 -53 64 -23
<< pdiffusion >>
rect 26 135 28 183
rect 35 135 37 183
rect 53 135 55 183
rect 62 135 64 183
<< pohmic >>
rect 0 -84 6 -77
rect 22 -84 34 -77
rect 50 -84 62 -77
rect 78 -84 99 -77
rect 0 -87 99 -84
<< nohmic >>
rect 0 214 99 217
rect 0 207 6 214
rect 22 207 34 214
rect 50 207 62 214
rect 78 207 99 214
<< ntransistor >>
rect 28 -53 35 -23
rect 55 -53 62 -23
<< ptransistor >>
rect 28 135 35 183
rect 55 135 62 183
<< polycontact >>
rect 45 49 61 65
rect 24 -13 40 3
<< ndiffcontact >>
rect 10 -53 26 -23
rect 64 -53 80 -23
<< pdiffcontact >>
rect 10 135 26 183
rect 37 135 53 183
rect 64 135 80 183
<< psubstratetap >>
rect 6 -84 22 -68
rect 34 -84 50 -68
rect 62 -84 78 -68
<< nsubstratetap >>
rect 6 198 22 214
rect 34 198 50 214
rect 62 198 78 214
<< metal1 >>
rect 0 214 99 217
rect 0 198 6 214
rect 22 198 34 214
rect 50 198 62 214
rect 78 198 99 214
rect 0 193 99 198
rect 10 183 26 193
rect 64 183 80 193
rect 37 85 47 135
rect 37 75 71 85
rect 71 39 81 71
rect 70 29 81 39
rect 70 -23 80 29
rect 10 -63 26 -53
rect 0 -68 99 -63
rect 0 -84 6 -68
rect 22 -84 34 -68
rect 50 -84 62 -68
rect 78 -84 99 -68
rect 0 -87 99 -84
<< m2contact >>
rect 71 71 85 85
rect 46 35 60 49
rect 24 3 38 17
<< metal2 >>
rect 24 194 36 221
rect 23 183 36 194
rect 24 135 37 183
rect 24 17 36 135
rect 48 65 60 221
rect 72 85 84 221
rect 48 49 61 65
rect 24 -13 38 3
rect 24 -68 36 -13
rect 23 -84 36 -68
rect 24 -91 36 -84
rect 48 -91 60 35
rect 72 -68 84 71
rect 71 -84 84 -68
rect 72 -91 84 -84
<< labels >>
rlabel metal1 99 193 99 217 7 Vdd!
rlabel metal1 0 193 0 217 3 Vdd!
rlabel metal2 24 221 36 221 5 A
rlabel metal2 48 221 60 221 5 B
rlabel metal2 72 221 84 221 5 Y
rlabel metal2 72 -91 84 -91 1 Y
rlabel metal2 48 -91 60 -91 1 B
rlabel metal2 24 -91 36 -91 1 A
rlabel metal1 0 -87 0 -63 3 GND!
rlabel metal1 99 -87 99 -63 7 GND!
<< end >>
