magic
tech c035u
timestamp 1385633360
<< nwell >>
rect 0 402 415 746
<< polysilicon >>
rect 63 691 70 719
rect 93 691 100 719
rect 144 704 211 711
rect 30 610 37 621
rect 30 388 37 562
rect 63 486 70 643
rect 93 612 100 643
rect 146 612 153 623
rect 187 612 194 645
rect 204 624 211 704
rect 249 691 256 719
rect 307 691 314 719
rect 249 624 256 643
rect 204 617 256 624
rect 249 612 256 617
rect 93 486 100 564
rect 146 486 153 564
rect 187 486 194 564
rect 249 486 256 564
rect 307 532 314 643
rect 375 612 382 675
rect 30 220 37 372
rect 63 331 70 438
rect 93 402 100 438
rect 146 428 153 438
rect 162 412 174 419
rect 93 395 134 402
rect 127 366 134 395
rect 167 366 174 412
rect 187 410 194 438
rect 249 428 256 438
rect 187 403 215 410
rect 208 366 215 403
rect 249 366 256 412
rect 63 288 70 315
rect 127 288 134 328
rect 30 182 37 190
rect 63 161 70 258
rect 127 220 134 258
rect 167 220 174 328
rect 208 220 215 328
rect 249 255 256 328
rect 249 248 263 255
rect 249 225 263 232
rect 249 220 256 225
rect 307 220 314 516
rect 339 486 346 539
rect 339 366 346 438
rect 339 288 346 328
rect 63 110 70 131
rect 127 127 134 190
rect 167 128 174 190
rect 208 161 215 190
rect 249 161 256 190
rect 307 180 314 190
rect 307 142 314 150
rect 339 142 346 258
rect 375 227 382 564
rect 365 220 382 227
rect 372 190 379 195
rect 365 188 379 190
rect 372 180 379 188
rect 372 142 379 150
rect 208 120 215 131
rect 249 120 256 131
<< ndiffusion >>
rect 122 328 127 366
rect 134 328 167 366
rect 174 328 181 366
rect 197 328 208 366
rect 215 328 249 366
rect 256 328 261 366
rect 58 258 63 288
rect 70 258 127 288
rect 134 258 145 288
rect 28 190 30 220
rect 37 190 42 220
rect 337 258 339 288
rect 346 258 352 288
rect 125 190 127 220
rect 134 190 167 220
rect 174 190 177 220
rect 241 190 249 220
rect 256 190 307 220
rect 314 190 318 220
rect 58 131 63 161
rect 70 131 75 161
rect 206 131 208 161
rect 215 131 249 161
rect 256 131 260 161
rect 369 150 372 180
rect 379 150 382 180
<< pdiffusion >>
rect 61 643 63 691
rect 70 643 72 691
rect 88 643 93 691
rect 100 643 102 691
rect 27 562 30 610
rect 37 562 42 610
rect 232 643 249 691
rect 256 643 266 691
rect 282 643 307 691
rect 314 643 317 691
rect 91 564 93 612
rect 100 564 128 612
rect 144 564 146 612
rect 153 564 163 612
rect 179 564 187 612
rect 194 564 196 612
rect 212 564 249 612
rect 256 564 258 612
rect 372 564 375 612
rect 382 564 392 612
rect 61 438 63 486
rect 70 438 73 486
rect 89 438 93 486
rect 100 438 102 486
rect 122 438 146 486
rect 153 438 161 486
rect 179 438 187 486
rect 194 438 196 486
rect 212 438 249 486
rect 256 438 259 486
rect 336 438 339 486
rect 346 438 352 486
<< ntransistor >>
rect 127 328 134 366
rect 167 328 174 366
rect 208 328 215 366
rect 249 328 256 366
rect 63 258 70 288
rect 127 258 134 288
rect 30 190 37 220
rect 339 258 346 288
rect 127 190 134 220
rect 167 190 174 220
rect 249 190 256 220
rect 307 190 314 220
rect 63 131 70 161
rect 208 131 215 161
rect 249 131 256 161
rect 372 150 379 180
<< ptransistor >>
rect 63 643 70 691
rect 93 643 100 691
rect 30 562 37 610
rect 249 643 256 691
rect 307 643 314 691
rect 93 564 100 612
rect 146 564 153 612
rect 187 564 194 612
rect 249 564 256 612
rect 375 564 382 612
rect 63 438 70 486
rect 93 438 100 486
rect 146 438 153 486
rect 187 438 194 486
rect 249 438 256 486
rect 339 438 346 486
<< polycontact >>
rect 128 695 144 711
rect 178 645 194 661
rect 366 675 382 691
rect 330 539 346 555
rect 302 516 318 532
rect 21 372 37 388
rect 146 412 162 428
rect 249 412 265 428
rect 59 315 75 331
rect 251 232 267 248
rect 330 328 346 366
rect 199 190 215 220
rect 307 150 323 180
rect 356 190 372 220
rect 122 111 138 127
rect 163 111 180 128
<< ndiffcontact >>
rect 106 328 122 366
rect 181 328 197 366
rect 261 328 277 366
rect 42 258 58 288
rect 145 258 161 288
rect 12 190 28 220
rect 42 190 58 220
rect 321 258 337 288
rect 352 258 368 288
rect 109 190 125 220
rect 177 190 193 220
rect 225 190 241 220
rect 318 190 334 220
rect 42 131 58 161
rect 75 131 91 161
rect 190 131 206 161
rect 260 131 276 161
rect 353 150 369 180
rect 382 150 398 180
<< pdiffcontact >>
rect 45 643 61 691
rect 72 643 88 691
rect 102 643 118 691
rect 11 562 27 610
rect 42 562 58 610
rect 216 643 232 691
rect 266 643 282 691
rect 317 643 333 691
rect 75 564 91 612
rect 128 564 144 612
rect 163 564 179 612
rect 196 564 212 612
rect 258 564 274 612
rect 356 564 372 612
rect 392 564 408 612
rect 45 438 61 486
rect 73 438 89 486
rect 102 438 122 486
rect 161 438 179 486
rect 196 438 212 486
rect 259 438 275 486
rect 320 438 336 486
rect 352 438 369 486
<< psubstratetap >>
rect 216 80 233 97
<< nsubstratetap >>
rect 226 727 243 744
<< metal1 >>
rect 0 782 415 792
rect 0 759 305 769
rect 321 759 415 769
rect 0 744 415 746
rect 0 727 226 744
rect 243 727 415 744
rect 0 721 415 727
rect 11 634 27 721
rect 45 691 61 721
rect 72 701 128 711
rect 72 691 88 701
rect 266 701 366 711
rect 266 691 282 701
rect 366 691 382 695
rect 11 633 28 634
rect 102 633 118 643
rect 11 621 118 633
rect 128 645 178 655
rect 11 610 27 621
rect 75 612 91 621
rect 11 511 27 562
rect 128 612 144 645
rect 216 633 232 643
rect 317 633 333 643
rect 392 633 408 721
rect 163 623 408 633
rect 163 612 179 623
rect 258 612 274 623
rect 392 612 408 623
rect 42 549 58 562
rect 128 549 144 564
rect 42 539 144 549
rect 196 554 212 564
rect 196 544 330 554
rect 102 516 276 526
rect 292 516 302 526
rect 356 526 372 564
rect 318 516 372 526
rect 11 501 89 511
rect 73 486 89 501
rect 102 486 122 516
rect 392 506 408 564
rect 161 496 275 506
rect 161 486 179 496
rect 259 486 275 496
rect 320 496 408 506
rect 320 486 336 496
rect 275 438 320 486
rect 45 428 61 438
rect 196 428 212 438
rect 352 428 369 438
rect 45 418 146 428
rect 162 418 212 428
rect 265 418 369 428
rect 60 390 197 402
rect 0 375 21 385
rect 60 353 73 390
rect 181 366 197 390
rect 12 341 73 353
rect 12 288 28 341
rect 59 314 75 315
rect 277 328 330 366
rect 106 318 122 328
rect 106 308 398 318
rect 12 258 42 288
rect 161 278 321 288
rect 12 220 28 258
rect 42 247 58 258
rect 352 248 368 258
rect 42 235 241 247
rect 225 220 241 235
rect 267 232 368 248
rect 58 190 109 220
rect 193 190 199 220
rect 334 190 356 220
rect 12 161 28 190
rect 382 180 398 308
rect 12 131 42 161
rect 91 151 190 161
rect 323 150 353 180
rect 12 101 30 131
rect 121 111 122 127
rect 260 121 276 131
rect 180 111 276 121
rect 0 97 415 101
rect 0 80 216 97
rect 233 80 415 97
rect 0 76 415 80
rect 0 53 59 63
rect 75 53 415 63
rect 0 30 415 40
rect 0 7 105 17
rect 121 7 415 17
<< m2contact >>
rect 305 756 321 772
rect 366 695 382 711
rect 276 516 292 532
rect 59 298 75 314
rect 105 111 121 127
rect 59 50 75 66
rect 105 3 121 19
<< metal2 >>
rect 278 532 290 799
rect 307 772 319 799
rect 307 711 319 756
rect 307 695 366 711
rect 59 66 75 298
rect 105 19 121 111
rect 278 0 290 516
rect 307 0 319 695
<< labels >>
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 1 Clock
rlabel metal1 0 7 0 17 1 nReset
rlabel metal1 415 7 415 17 7 nReset
rlabel metal1 415 30 415 40 7 Test
rlabel metal1 415 53 415 63 7 Clock
rlabel metal1 415 76 415 101 7 GND!
rlabel metal2 307 0 319 0 1 Q
rlabel metal2 278 0 290 0 1 nQ
rlabel metal1 415 759 415 769 7 Q
rlabel metal1 415 782 415 792 7 ScanReturn
rlabel metal2 307 799 319 799 5 Q
rlabel metal2 278 799 290 799 5 nQ
rlabel metal1 0 759 0 769 3 Q
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 375 0 385 3 D
<< end >>
