magic
tech c035u
timestamp 1385637965
<< nwell >>
rect 0 402 180 746
<< polysilicon >>
rect 115 618 122 627
rect 63 539 70 547
rect 83 539 90 549
rect 63 481 70 491
rect 33 460 40 468
rect 33 391 40 412
rect 33 365 40 375
rect 33 327 40 335
rect 63 330 70 465
rect 63 304 70 314
rect 83 304 90 491
rect 115 481 122 570
rect 63 266 70 274
rect 83 264 90 274
rect 115 243 122 465
rect 115 205 122 213
<< ndiffusion >>
rect 31 335 33 365
rect 40 335 42 365
rect 61 274 63 304
rect 70 274 83 304
rect 90 274 92 304
rect 113 213 115 243
rect 122 213 124 243
<< pdiffusion >>
rect 113 570 115 618
rect 122 570 124 618
rect 61 491 63 539
rect 70 491 83 539
rect 90 491 92 539
rect 31 412 33 460
rect 40 412 42 460
<< ntransistor >>
rect 33 335 40 365
rect 63 274 70 304
rect 83 274 90 304
rect 115 213 122 243
<< ptransistor >>
rect 115 570 122 618
rect 63 491 70 539
rect 83 491 90 539
rect 33 412 40 460
<< polycontact >>
rect 83 549 99 565
rect 57 465 73 481
rect 32 375 48 391
rect 57 314 73 330
rect 115 465 131 481
rect 83 248 99 264
<< ndiffcontact >>
rect 15 335 31 365
rect 42 335 58 365
rect 45 274 61 304
rect 92 274 108 304
rect 97 213 113 243
rect 124 213 140 243
<< pdiffcontact >>
rect 96 570 113 618
rect 124 570 141 618
rect 45 491 61 539
rect 92 491 108 539
rect 15 412 31 460
rect 42 412 58 460
<< metal1 >>
rect 0 782 180 792
rect 0 759 180 769
rect 0 721 180 746
rect 15 460 31 721
rect 45 539 61 721
rect 124 618 141 721
rect 83 570 96 618
rect 83 565 99 570
rect 42 465 57 481
rect 42 460 58 465
rect 92 425 105 491
rect 115 464 131 465
rect 92 408 149 425
rect 31 375 32 391
rect 15 101 31 335
rect 42 330 58 335
rect 42 314 57 330
rect 92 304 105 408
rect 45 101 61 274
rect 83 243 99 248
rect 83 213 97 243
rect 124 101 140 213
rect 0 76 180 101
rect 0 53 180 63
rect 0 30 180 40
rect 0 7 180 17
<< m2contact >>
rect 115 448 131 464
rect 149 408 165 425
rect 15 375 31 391
<< metal2 >>
rect 15 391 31 799
rect 15 0 31 375
rect 79 464 95 799
rect 79 448 115 464
rect 79 0 95 448
rect 149 425 165 799
rect 149 0 165 408
<< labels >>
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 180 7 180 17 8 nReset
rlabel metal1 180 30 180 40 7 Test
rlabel metal1 180 53 180 63 7 Clock
rlabel metal1 180 76 180 101 7 GND!
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 180 782 180 792 6 ScanReturn
rlabel metal1 180 759 180 769 7 Scan
rlabel metal1 180 721 180 746 7 Vdd!
rlabel metal2 149 0 165 0 1 Y
rlabel metal2 15 0 31 0 1 A
rlabel metal2 79 0 95 0 1 Enable
rlabel metal2 149 799 165 799 5 Y
rlabel metal2 15 799 31 799 5 A
rlabel metal2 79 799 95 799 5 Enable
<< end >>
