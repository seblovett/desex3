magic
tech c035u
timestamp 1385918469
<< nwell >>
rect 0 402 264 746
<< polysilicon >>
rect 51 697 58 711
rect 24 669 31 677
rect 51 669 58 681
rect 147 669 154 677
rect 177 669 184 677
rect 232 669 239 677
rect 24 591 31 621
rect 51 591 58 621
rect 106 591 113 637
rect 24 249 31 543
rect 24 201 31 231
rect 51 201 58 543
rect 106 201 113 543
rect 147 533 154 621
rect 177 591 184 621
rect 232 561 239 621
rect 238 545 239 561
rect 147 227 154 517
rect 177 279 184 543
rect 24 141 31 171
rect 51 141 58 171
rect 106 161 113 171
rect 147 141 154 211
rect 177 201 184 263
rect 232 217 239 545
rect 177 141 184 171
rect 232 141 239 201
rect 24 103 31 111
rect 51 103 58 111
rect 147 103 154 111
rect 177 103 184 111
rect 232 103 239 111
<< ndiffusion >>
rect 22 171 24 201
rect 31 171 51 201
rect 58 171 60 201
rect 104 171 106 201
rect 113 171 115 201
rect 175 171 177 201
rect 184 171 186 201
rect 22 111 24 141
rect 31 111 33 141
rect 49 111 51 141
rect 58 111 60 141
rect 145 111 147 141
rect 154 111 177 141
rect 184 111 186 141
rect 230 111 232 141
rect 239 111 241 141
<< pdiffusion >>
rect 22 621 24 669
rect 31 621 51 669
rect 58 621 60 669
rect 145 621 147 669
rect 154 621 159 669
rect 175 621 177 669
rect 184 621 186 669
rect 202 621 232 669
rect 239 621 241 669
rect 22 543 24 591
rect 31 543 33 591
rect 49 543 51 591
rect 58 543 60 591
rect 76 543 106 591
rect 113 543 115 591
rect 175 543 177 591
rect 184 543 186 591
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 174 86
rect 190 76 202 86
rect 218 76 230 86
rect 246 76 264 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
rect 50 736 62 746
rect 78 736 90 746
rect 106 736 118 746
rect 134 736 146 746
rect 162 736 174 746
rect 190 736 202 746
rect 218 736 230 746
rect 246 736 264 746
<< ntransistor >>
rect 24 171 31 201
rect 51 171 58 201
rect 106 171 113 201
rect 177 171 184 201
rect 24 111 31 141
rect 51 111 58 141
rect 147 111 154 141
rect 177 111 184 141
rect 232 111 239 141
<< ptransistor >>
rect 24 621 31 669
rect 51 621 58 669
rect 147 621 154 669
rect 177 621 184 669
rect 232 621 239 669
rect 24 543 31 591
rect 51 543 58 591
rect 106 543 113 591
rect 177 543 184 591
<< polycontact >>
rect 47 681 63 697
rect 101 637 117 653
rect 22 231 40 249
rect 222 545 238 561
rect 138 517 154 533
rect 168 263 184 279
rect 138 211 154 227
rect 101 145 117 161
rect 223 201 239 217
<< ndiffcontact >>
rect 6 171 22 201
rect 60 171 76 201
rect 88 171 104 201
rect 115 171 131 201
rect 159 171 175 201
rect 186 171 202 201
rect 6 111 22 141
rect 33 111 49 141
rect 60 111 76 141
rect 129 111 145 141
rect 186 111 202 141
rect 214 111 230 141
rect 241 111 257 141
<< pdiffcontact >>
rect 6 621 22 669
rect 60 621 76 669
rect 129 621 145 669
rect 159 621 175 669
rect 186 621 202 669
rect 241 621 257 669
rect 6 543 22 591
rect 33 543 49 591
rect 60 543 76 591
rect 115 543 131 591
rect 159 543 175 591
rect 186 543 202 591
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
rect 174 76 190 92
rect 202 76 218 92
rect 230 76 246 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
rect 62 730 78 746
rect 90 730 106 746
rect 118 730 134 746
rect 146 730 162 746
rect 174 730 190 746
rect 202 730 218 746
rect 230 730 246 746
<< metal1 >>
rect 0 782 264 792
rect 0 759 264 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 62 746
rect 78 730 90 746
rect 106 730 118 746
rect 134 730 146 746
rect 162 730 174 746
rect 190 730 202 746
rect 218 730 230 746
rect 246 730 264 746
rect 0 721 264 730
rect 9 669 19 721
rect 132 669 142 721
rect 189 669 199 721
rect 76 640 101 650
rect 9 611 19 621
rect 135 611 145 621
rect 162 611 172 621
rect 9 601 73 611
rect 135 601 152 611
rect 162 601 231 611
rect 9 591 19 601
rect 63 591 73 601
rect 142 591 152 601
rect 142 581 159 591
rect 221 561 231 601
rect 243 585 253 621
rect 221 545 222 561
rect 36 276 46 543
rect 118 530 128 543
rect 192 533 202 543
rect 118 519 138 530
rect 36 266 168 276
rect 63 201 73 266
rect 91 217 138 227
rect 91 201 101 217
rect 192 201 202 227
rect 131 181 159 191
rect 9 141 19 171
rect 36 151 101 161
rect 36 141 46 151
rect 131 141 141 181
rect 222 201 223 217
rect 222 161 232 201
rect 189 151 232 161
rect 189 141 199 151
rect 244 141 254 177
rect 9 101 19 111
rect 63 101 73 111
rect 132 101 142 111
rect 217 101 227 111
rect 0 92 264 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 174 92
rect 190 76 202 92
rect 218 76 230 92
rect 246 76 264 92
rect 0 53 264 63
rect 0 30 264 40
rect 0 7 264 17
<< m2contact >>
rect 47 697 61 711
rect 241 571 255 585
rect 191 519 205 533
rect 24 217 38 231
rect 191 227 205 241
rect 242 177 256 191
<< metal2 >>
rect 24 231 36 799
rect 48 711 60 799
rect 24 0 36 217
rect 48 0 60 697
rect 192 533 204 799
rect 240 585 252 799
rect 240 571 241 585
rect 192 241 204 519
rect 192 0 204 227
rect 240 191 252 571
rect 240 177 242 191
rect 240 0 252 177
<< labels >>
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 264 76 264 101 7 GND!
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 264 53 264 63 7 Clock
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 264 30 264 40 7 Test
rlabel metal2 24 0 36 0 1 A
rlabel metal2 48 0 60 0 1 B
rlabel metal2 192 0 204 0 1 C
rlabel metal2 240 0 252 0 1 S
rlabel metal1 0 7 0 17 3 nReset
rlabel metal1 264 7 264 17 7 nReset
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 264 721 264 746 7 Vdd!
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 264 759 264 769 7 Scan
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 264 782 264 792 7 ScanReturn
rlabel metal2 240 799 252 799 5 S
rlabel metal2 192 799 204 799 5 C
rlabel metal2 48 799 60 799 5 B
rlabel metal2 24 799 36 799 5 A
<< end >>
