magic
tech c035u
timestamp 1385930293
<< nwell >>
rect 202 392 1464 736
rect 405 391 451 392
rect 742 391 788 392
rect 1079 391 1125 392
<< polysilicon >>
rect 538 682 545 690
rect 565 682 572 690
rect 592 682 599 690
rect 619 682 626 690
rect 875 682 882 690
rect 902 682 909 690
rect 929 682 936 690
rect 956 682 963 690
rect 1212 682 1219 690
rect 1239 682 1246 690
rect 1266 682 1273 690
rect 1293 682 1300 690
rect 480 604 487 612
rect 507 604 514 612
rect 425 549 432 557
rect 370 450 377 458
rect 817 604 824 612
rect 844 604 851 612
rect 762 549 769 557
rect 707 450 714 458
rect 1154 604 1161 612
rect 1181 604 1188 612
rect 1099 549 1106 557
rect 1044 450 1051 458
rect 1394 506 1396 522
rect 1389 461 1396 506
rect 370 378 377 392
rect 425 378 432 392
rect 480 379 487 392
rect 375 362 377 378
rect 430 362 432 378
rect 485 375 487 379
rect 507 375 514 392
rect 538 379 545 392
rect 485 368 514 375
rect 485 363 487 368
rect 543 375 545 379
rect 565 375 572 392
rect 592 375 599 392
rect 619 375 626 392
rect 707 378 714 392
rect 762 378 769 392
rect 817 379 824 392
rect 543 368 626 375
rect 543 363 545 368
rect 370 301 377 362
rect 425 301 432 362
rect 480 301 487 363
rect 538 301 545 363
rect 565 301 572 368
rect 712 362 714 378
rect 767 362 769 378
rect 822 375 824 379
rect 844 375 851 392
rect 875 379 882 392
rect 822 368 851 375
rect 822 363 824 368
rect 880 375 882 379
rect 902 375 909 392
rect 929 375 936 392
rect 956 375 963 392
rect 1044 378 1051 392
rect 1099 378 1106 392
rect 1154 379 1161 392
rect 880 368 963 375
rect 880 363 882 368
rect 707 301 714 362
rect 762 301 769 362
rect 817 301 824 363
rect 875 301 882 363
rect 902 301 909 368
rect 1049 362 1051 378
rect 1104 362 1106 378
rect 1159 375 1161 379
rect 1181 375 1188 392
rect 1212 379 1219 392
rect 1159 368 1188 375
rect 1159 363 1161 368
rect 1217 375 1219 379
rect 1239 375 1246 392
rect 1266 375 1273 392
rect 1293 375 1300 392
rect 1217 368 1300 375
rect 1217 363 1219 368
rect 1044 301 1051 362
rect 1099 301 1106 362
rect 1154 301 1161 363
rect 1212 301 1219 363
rect 1239 301 1246 368
rect 1389 309 1396 413
rect 370 273 377 281
rect 425 239 432 247
rect 480 147 487 155
rect 707 273 714 281
rect 762 239 769 247
rect 817 147 824 155
rect 1044 273 1051 281
rect 1099 239 1106 247
rect 1154 147 1161 155
rect 1389 271 1396 279
rect 538 93 545 101
rect 565 93 572 101
rect 875 93 882 101
rect 902 93 909 101
rect 1212 93 1219 101
rect 1239 93 1246 101
<< ndiffusion >>
rect 368 281 370 301
rect 377 281 379 301
rect 423 247 425 301
rect 432 247 434 301
rect 478 155 480 301
rect 487 155 489 301
rect 536 101 538 301
rect 545 101 547 301
rect 563 101 565 301
rect 572 101 574 301
rect 705 281 707 301
rect 714 281 716 301
rect 760 247 762 301
rect 769 247 771 301
rect 815 155 817 301
rect 824 155 826 301
rect 873 101 875 301
rect 882 101 884 301
rect 900 101 902 301
rect 909 101 911 301
rect 1042 281 1044 301
rect 1051 281 1053 301
rect 1097 247 1099 301
rect 1106 247 1108 301
rect 1152 155 1154 301
rect 1161 155 1163 301
rect 1210 101 1212 301
rect 1219 101 1221 301
rect 1237 101 1239 301
rect 1246 101 1248 301
rect 1387 279 1389 309
rect 1396 279 1398 309
<< pdiffusion >>
rect 368 392 370 450
rect 377 392 379 450
rect 423 392 425 549
rect 432 392 434 549
rect 478 392 480 604
rect 487 392 489 604
rect 505 392 507 604
rect 514 392 516 604
rect 536 392 538 682
rect 545 392 547 682
rect 563 392 565 682
rect 572 392 574 682
rect 590 392 592 682
rect 599 392 601 682
rect 617 392 619 682
rect 626 392 628 682
rect 705 392 707 450
rect 714 392 716 450
rect 760 392 762 549
rect 769 392 771 549
rect 815 392 817 604
rect 824 392 826 604
rect 842 392 844 604
rect 851 392 853 604
rect 873 392 875 682
rect 882 392 884 682
rect 900 392 902 682
rect 909 392 911 682
rect 927 392 929 682
rect 936 392 938 682
rect 954 392 956 682
rect 963 392 965 682
rect 1042 392 1044 450
rect 1051 392 1053 450
rect 1097 392 1099 549
rect 1106 392 1108 549
rect 1152 392 1154 604
rect 1161 392 1163 604
rect 1179 392 1181 604
rect 1188 392 1190 604
rect 1210 392 1212 682
rect 1219 392 1221 682
rect 1237 392 1239 682
rect 1246 392 1248 682
rect 1264 392 1266 682
rect 1273 392 1275 682
rect 1291 392 1293 682
rect 1300 392 1302 682
rect 1387 413 1389 461
rect 1396 413 1398 461
<< pohmic >>
rect 320 66 326 76
rect 342 66 354 76
rect 370 66 382 76
rect 398 66 410 76
rect 426 66 438 76
rect 454 66 466 76
rect 482 66 494 76
rect 510 66 522 76
rect 538 66 550 76
rect 567 66 579 76
rect 595 66 607 76
rect 623 66 635 76
rect 651 66 663 76
rect 679 66 691 76
rect 707 66 719 76
rect 735 66 747 76
rect 763 66 775 76
rect 791 66 803 76
rect 819 66 831 76
rect 847 66 859 76
rect 875 66 887 76
rect 904 66 916 76
rect 932 66 944 76
rect 960 66 972 76
rect 988 66 1000 76
rect 1016 66 1028 76
rect 1044 66 1056 76
rect 1072 66 1084 76
rect 1100 66 1112 76
rect 1128 66 1140 76
rect 1156 66 1168 76
rect 1184 66 1196 76
rect 1212 66 1224 76
rect 1241 66 1253 76
rect 1269 66 1281 76
rect 1297 66 1309 76
rect 1325 66 1337 76
rect 1353 66 1365 76
rect 1381 66 1393 76
rect 1409 66 1421 76
rect 1437 66 1464 76
<< nohmic >>
rect 202 726 214 736
rect 230 726 242 736
rect 258 726 270 736
rect 286 726 298 736
rect 314 726 326 736
rect 342 726 354 736
rect 370 726 382 736
rect 398 726 410 736
rect 426 726 438 736
rect 454 726 466 736
rect 482 726 494 736
rect 510 726 522 736
rect 538 726 550 736
rect 567 726 579 736
rect 595 726 607 736
rect 623 726 635 736
rect 651 726 663 736
rect 679 726 691 736
rect 707 726 719 736
rect 735 726 747 736
rect 763 726 775 736
rect 791 726 803 736
rect 819 726 831 736
rect 847 726 859 736
rect 875 726 887 736
rect 904 726 916 736
rect 932 726 944 736
rect 960 726 972 736
rect 988 726 1000 736
rect 1016 726 1028 736
rect 1044 726 1056 736
rect 1072 726 1084 736
rect 1100 726 1112 736
rect 1128 726 1140 736
rect 1156 726 1168 736
rect 1184 726 1196 736
rect 1212 726 1224 736
rect 1241 726 1253 736
rect 1269 726 1281 736
rect 1297 726 1309 736
rect 1325 726 1337 736
rect 1353 726 1365 736
rect 1381 726 1393 736
rect 1409 726 1421 736
rect 1437 726 1464 736
<< ntransistor >>
rect 370 281 377 301
rect 425 247 432 301
rect 480 155 487 301
rect 538 101 545 301
rect 565 101 572 301
rect 707 281 714 301
rect 762 247 769 301
rect 817 155 824 301
rect 875 101 882 301
rect 902 101 909 301
rect 1044 281 1051 301
rect 1099 247 1106 301
rect 1154 155 1161 301
rect 1212 101 1219 301
rect 1239 101 1246 301
rect 1389 279 1396 309
<< ptransistor >>
rect 370 392 377 450
rect 425 392 432 549
rect 480 392 487 604
rect 507 392 514 604
rect 538 392 545 682
rect 565 392 572 682
rect 592 392 599 682
rect 619 392 626 682
rect 707 392 714 450
rect 762 392 769 549
rect 817 392 824 604
rect 844 392 851 604
rect 875 392 882 682
rect 902 392 909 682
rect 929 392 936 682
rect 956 392 963 682
rect 1044 392 1051 450
rect 1099 392 1106 549
rect 1154 392 1161 604
rect 1181 392 1188 604
rect 1212 392 1219 682
rect 1239 392 1246 682
rect 1266 392 1273 682
rect 1293 392 1300 682
rect 1389 413 1396 461
<< polycontact >>
rect 1378 506 1394 522
rect 359 362 375 378
rect 414 362 430 378
rect 469 363 485 379
rect 527 363 543 379
rect 696 362 712 378
rect 751 362 767 378
rect 806 363 822 379
rect 864 363 880 379
rect 1033 362 1049 378
rect 1088 362 1104 378
rect 1143 363 1159 379
rect 1201 363 1217 379
<< ndiffcontact >>
rect 352 281 368 301
rect 379 281 395 301
rect 407 247 423 301
rect 434 247 450 301
rect 462 155 478 301
rect 489 155 505 301
rect 520 101 536 301
rect 547 101 563 301
rect 574 101 590 301
rect 689 281 705 301
rect 716 281 732 301
rect 744 247 760 301
rect 771 247 787 301
rect 799 155 815 301
rect 826 155 842 301
rect 857 101 873 301
rect 884 101 900 301
rect 911 101 927 301
rect 1026 281 1042 301
rect 1053 281 1069 301
rect 1081 247 1097 301
rect 1108 247 1124 301
rect 1136 155 1152 301
rect 1163 155 1179 301
rect 1194 101 1210 301
rect 1221 101 1237 301
rect 1248 101 1264 301
rect 1371 279 1387 309
rect 1398 279 1414 309
<< pdiffcontact >>
rect 519 604 536 682
rect 352 392 368 450
rect 379 392 395 450
rect 407 392 423 549
rect 434 392 450 549
rect 462 392 478 604
rect 489 392 505 604
rect 516 392 536 604
rect 547 392 563 682
rect 574 392 590 682
rect 601 392 617 682
rect 628 392 644 682
rect 856 604 873 682
rect 689 392 705 450
rect 716 392 732 450
rect 744 392 760 549
rect 771 392 787 549
rect 799 392 815 604
rect 826 392 842 604
rect 853 392 873 604
rect 884 392 900 682
rect 911 392 927 682
rect 938 392 954 682
rect 965 392 981 682
rect 1193 604 1210 682
rect 1026 392 1042 450
rect 1053 392 1069 450
rect 1081 392 1097 549
rect 1108 392 1124 549
rect 1136 392 1152 604
rect 1163 392 1179 604
rect 1190 392 1210 604
rect 1221 392 1237 682
rect 1248 392 1264 682
rect 1275 392 1291 682
rect 1302 392 1318 682
rect 1371 413 1387 461
rect 1398 413 1414 461
<< psubstratetap >>
rect 326 66 342 82
rect 354 66 370 82
rect 382 66 398 82
rect 410 66 426 82
rect 438 66 454 82
rect 466 66 482 82
rect 494 66 510 82
rect 522 66 538 82
rect 550 66 567 82
rect 579 66 595 82
rect 607 66 623 82
rect 635 66 651 82
rect 663 66 679 82
rect 691 66 707 82
rect 719 66 735 82
rect 747 66 763 82
rect 775 66 791 82
rect 803 66 819 82
rect 831 66 847 82
rect 859 66 875 82
rect 887 66 904 82
rect 916 66 932 82
rect 944 66 960 82
rect 972 66 988 82
rect 1000 66 1016 82
rect 1028 66 1044 82
rect 1056 66 1072 82
rect 1084 66 1100 82
rect 1112 66 1128 82
rect 1140 66 1156 82
rect 1168 66 1184 82
rect 1196 66 1212 82
rect 1224 66 1241 82
rect 1253 66 1269 82
rect 1281 66 1297 82
rect 1309 66 1325 82
rect 1337 66 1353 82
rect 1365 66 1381 82
rect 1393 66 1409 82
rect 1421 66 1437 82
<< nsubstratetap >>
rect 214 720 230 736
rect 242 720 258 736
rect 270 720 286 736
rect 298 720 314 736
rect 326 720 342 736
rect 354 720 370 736
rect 382 720 398 736
rect 410 720 426 736
rect 438 720 454 736
rect 466 720 482 736
rect 494 720 510 736
rect 522 720 538 736
rect 550 720 567 736
rect 579 720 595 736
rect 607 720 623 736
rect 635 720 651 736
rect 663 720 679 736
rect 691 720 707 736
rect 719 720 735 736
rect 747 720 763 736
rect 775 720 791 736
rect 803 720 819 736
rect 831 720 847 736
rect 859 720 875 736
rect 887 720 904 736
rect 916 720 932 736
rect 944 720 960 736
rect 972 720 988 736
rect 1000 720 1016 736
rect 1028 720 1044 736
rect 1056 720 1072 736
rect 1084 720 1100 736
rect 1112 720 1128 736
rect 1140 720 1156 736
rect 1168 720 1184 736
rect 1196 720 1212 736
rect 1224 720 1241 736
rect 1253 720 1269 736
rect 1281 720 1297 736
rect 1309 720 1325 736
rect 1337 720 1353 736
rect 1365 720 1381 736
rect 1393 720 1409 736
rect 1421 720 1437 736
<< metal1 >>
rect 229 772 1356 782
rect 1400 772 1464 782
rect 229 749 1464 759
rect 200 720 214 736
rect 230 720 242 736
rect 258 720 270 736
rect 286 720 298 736
rect 314 720 326 736
rect 342 720 354 736
rect 370 720 382 736
rect 398 720 410 736
rect 426 720 438 736
rect 454 720 466 736
rect 482 720 494 736
rect 510 720 522 736
rect 538 720 550 736
rect 567 720 579 736
rect 595 720 607 736
rect 623 720 635 736
rect 651 720 663 736
rect 679 720 691 736
rect 707 720 719 736
rect 735 720 747 736
rect 763 720 775 736
rect 791 720 803 736
rect 819 720 831 736
rect 847 720 859 736
rect 875 720 887 736
rect 904 720 916 736
rect 932 720 944 736
rect 960 720 972 736
rect 988 720 1000 736
rect 1016 720 1028 736
rect 1044 720 1056 736
rect 1072 720 1084 736
rect 1100 720 1112 736
rect 1128 720 1140 736
rect 1156 720 1168 736
rect 1184 720 1196 736
rect 1212 720 1224 736
rect 1241 720 1253 736
rect 1269 720 1281 736
rect 1297 720 1309 736
rect 1325 720 1337 736
rect 1353 720 1365 736
rect 1381 720 1393 736
rect 1409 720 1421 736
rect 1437 720 1464 736
rect 200 711 1464 720
rect 352 450 368 711
rect 407 549 423 711
rect 462 604 478 711
rect 516 682 536 711
rect 574 682 590 711
rect 628 682 644 711
rect 516 604 519 682
rect 689 450 705 711
rect 744 549 760 711
rect 799 604 815 711
rect 853 682 873 711
rect 911 682 927 711
rect 965 682 981 711
rect 853 604 856 682
rect 1026 450 1042 711
rect 1081 549 1097 711
rect 1136 604 1152 711
rect 1190 682 1210 711
rect 1248 682 1264 711
rect 1302 682 1318 711
rect 1190 604 1193 682
rect 1380 522 1394 528
rect 1404 461 1414 711
rect 277 365 359 375
rect 263 353 277 363
rect 385 375 395 392
rect 385 365 414 375
rect 385 301 395 365
rect 440 376 450 392
rect 440 366 469 376
rect 440 301 450 366
rect 495 376 505 392
rect 495 366 527 376
rect 495 301 505 366
rect 553 377 563 392
rect 607 379 617 392
rect 553 367 606 377
rect 553 301 563 367
rect 667 365 696 375
rect 722 375 732 392
rect 722 365 751 375
rect 722 301 732 365
rect 777 376 787 392
rect 777 366 806 376
rect 777 301 787 366
rect 832 376 842 392
rect 832 366 864 376
rect 832 301 842 366
rect 890 377 900 392
rect 944 379 954 392
rect 890 367 944 377
rect 890 301 900 367
rect 1022 365 1033 375
rect 1059 375 1069 392
rect 1059 365 1088 375
rect 1059 301 1069 365
rect 1114 376 1124 392
rect 1114 366 1143 376
rect 1114 301 1124 366
rect 1169 376 1179 392
rect 1169 366 1201 376
rect 1169 301 1179 366
rect 1227 377 1237 392
rect 1281 379 1291 392
rect 1227 367 1279 377
rect 1227 301 1237 367
rect 1371 309 1381 413
rect 352 91 368 281
rect 407 91 423 247
rect 462 91 478 155
rect 520 91 536 101
rect 574 91 590 101
rect 689 91 705 281
rect 744 91 760 247
rect 799 91 815 155
rect 857 91 873 101
rect 911 91 927 101
rect 1026 91 1042 281
rect 1081 91 1097 247
rect 1136 91 1152 155
rect 1194 91 1210 101
rect 1248 91 1264 101
rect 1398 91 1408 279
rect 320 82 1464 91
rect 320 66 326 82
rect 342 66 354 82
rect 370 66 382 82
rect 398 66 410 82
rect 426 66 438 82
rect 454 66 466 82
rect 482 66 494 82
rect 510 66 522 82
rect 538 66 550 82
rect 567 66 579 82
rect 595 66 607 82
rect 623 66 635 82
rect 651 66 663 82
rect 679 66 691 82
rect 707 66 719 82
rect 735 66 747 82
rect 763 66 775 82
rect 791 66 803 82
rect 819 66 831 82
rect 847 66 859 82
rect 875 66 887 82
rect 904 66 916 82
rect 932 66 944 82
rect 960 66 972 82
rect 988 66 1000 82
rect 1016 66 1028 82
rect 1044 66 1056 82
rect 1072 66 1084 82
rect 1100 66 1112 82
rect 1128 66 1140 82
rect 1156 66 1168 82
rect 1184 66 1196 82
rect 1212 66 1224 82
rect 1241 66 1253 82
rect 1269 66 1281 82
rect 1297 66 1309 82
rect 1325 66 1337 82
rect 1353 66 1365 82
rect 1381 66 1393 82
rect 1409 66 1421 82
rect 1437 66 1464 82
rect 239 33 253 43
rect 620 43 1464 53
rect 253 20 653 30
rect 959 20 1464 30
rect 301 -3 1009 7
rect 1294 -3 1304 7
rect 1318 -3 1464 7
<< m2contact >>
rect 215 770 229 784
rect 1356 771 1370 785
rect 1386 771 1400 785
rect 215 746 229 760
rect 0 711 200 736
rect 1380 528 1394 542
rect 1357 447 1371 461
rect 263 363 277 377
rect 263 339 277 353
rect 606 365 620 379
rect 653 363 667 377
rect 944 365 958 379
rect 1008 363 1022 377
rect 1279 365 1293 379
rect 239 43 253 57
rect 606 41 620 55
rect 239 19 253 33
rect 653 18 667 32
rect 945 19 959 33
rect 239 -5 253 9
rect 263 -5 277 9
rect 287 -5 301 9
rect 1009 -5 1023 9
rect 1280 -5 1294 9
rect 1304 -5 1318 9
<< metal2 >>
rect 0 736 200 789
rect 216 784 228 789
rect 0 -10 200 711
rect 216 -10 228 746
rect 240 57 252 789
rect 264 377 276 789
rect 264 353 276 363
rect 240 33 252 43
rect 240 9 252 19
rect 264 9 276 339
rect 288 9 300 789
rect 1358 461 1370 771
rect 1386 542 1398 771
rect 1394 528 1398 542
rect 607 55 619 365
rect 654 32 666 363
rect 946 33 958 365
rect 1010 9 1022 363
rect 1281 9 1293 365
rect 1294 -5 1304 9
rect 240 -10 252 -5
rect 264 -10 276 -5
rect 288 -10 300 -5
<< labels >>
rlabel metal2 0 789 200 789 5 Vdd!
rlabel metal2 0 -10 200 -10 1 Vdd!
rlabel metal1 1464 711 1464 736 7 Vdd!
rlabel metal1 1464 749 1464 759 7 SDI
rlabel metal1 1464 772 1464 782 7 nSDO
rlabel metal1 1464 43 1464 53 7 ClockOut
rlabel metal1 1464 20 1464 30 7 TestOut
rlabel metal1 1464 -3 1464 7 7 nResetOut
rlabel metal1 1464 66 1464 91 7 GND!
rlabel metal2 216 -10 228 -10 1 SDI
rlabel metal2 240 -10 252 -10 1 Test
rlabel metal2 264 -10 276 -10 1 Clock
rlabel metal2 288 -10 300 -10 1 nReset
rlabel metal2 288 789 300 789 5 nReset
rlabel metal2 240 789 252 789 5 Test
rlabel metal2 264 789 276 789 5 Clock
rlabel metal2 216 789 228 789 5 SDO
<< end >>
