magic
tech c035u
timestamp 1386235180
<< nwell >>
rect 0 401 288 799
<< pwell >>
rect 0 0 288 401
<< polysilicon >>
rect 216 681 221 697
rect 28 671 35 679
rect 58 671 65 679
rect 88 671 95 679
rect 132 671 139 679
rect 162 671 169 679
rect 189 671 196 679
rect 216 671 223 681
rect 28 375 35 623
rect 58 553 65 623
rect 88 539 95 623
rect 132 553 139 623
rect 88 523 93 539
rect 58 381 65 505
rect 28 235 35 359
rect 58 335 65 365
rect 88 335 95 523
rect 132 381 139 505
rect 162 381 169 623
rect 189 501 196 623
rect 132 335 139 365
rect 88 319 93 335
rect 58 235 65 305
rect 88 235 95 319
rect 132 235 139 305
rect 162 235 169 365
rect 189 355 196 485
rect 189 235 196 339
rect 216 235 223 623
rect 246 583 251 599
rect 246 553 253 583
rect 246 358 253 505
rect 246 275 253 328
rect 251 259 253 275
rect 28 197 35 205
rect 58 197 65 205
rect 88 197 95 205
rect 132 197 139 205
rect 162 197 169 205
rect 189 197 196 205
rect 216 197 223 205
<< ndiffusion >>
rect 56 305 58 335
rect 65 305 67 335
rect 130 305 132 335
rect 139 305 141 335
rect 244 328 246 358
rect 253 328 255 358
rect 26 205 28 235
rect 35 205 58 235
rect 65 205 67 235
rect 83 205 88 235
rect 95 205 114 235
rect 130 205 132 235
rect 139 205 162 235
rect 169 205 171 235
rect 187 205 189 235
rect 196 205 216 235
rect 223 205 225 235
<< pdiffusion >>
rect 26 623 28 671
rect 35 623 40 671
rect 56 623 58 671
rect 65 623 67 671
rect 83 623 88 671
rect 95 623 114 671
rect 130 623 132 671
rect 139 623 141 671
rect 157 623 162 671
rect 169 623 171 671
rect 187 623 189 671
rect 196 623 198 671
rect 214 623 216 671
rect 223 623 225 671
rect 56 505 58 553
rect 65 505 67 553
rect 130 505 132 553
rect 139 505 141 553
rect 244 505 246 553
rect 253 505 255 553
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 174 86
rect 190 79 202 86
rect 218 79 230 86
rect 246 79 258 86
rect 274 79 288 86
rect 0 76 288 79
<< nohmic >>
rect 0 743 288 746
rect 0 736 6 743
rect 22 736 34 743
rect 50 736 62 743
rect 78 736 90 743
rect 106 736 118 743
rect 134 736 146 743
rect 162 736 174 743
rect 190 736 202 743
rect 218 736 230 743
rect 246 736 258 743
rect 274 736 288 743
<< ntransistor >>
rect 58 305 65 335
rect 132 305 139 335
rect 246 328 253 358
rect 28 205 35 235
rect 58 205 65 235
rect 88 205 95 235
rect 132 205 139 235
rect 162 205 169 235
rect 189 205 196 235
rect 216 205 223 235
<< ptransistor >>
rect 28 623 35 671
rect 58 623 65 671
rect 88 623 95 671
rect 132 623 139 671
rect 162 623 169 671
rect 189 623 196 671
rect 216 623 223 671
rect 58 505 65 553
rect 132 505 139 553
rect 246 505 253 553
<< polycontact >>
rect 221 681 237 697
rect 93 523 109 539
rect 24 359 40 375
rect 54 365 70 381
rect 180 485 196 501
rect 127 365 143 381
rect 158 365 174 381
rect 93 319 109 335
rect 180 339 196 355
rect 251 583 267 599
rect 235 259 251 275
<< ndiffcontact >>
rect 40 305 56 335
rect 67 305 83 335
rect 114 305 130 335
rect 141 305 157 335
rect 228 328 244 358
rect 255 328 271 358
rect 10 205 26 235
rect 67 205 83 235
rect 114 205 130 235
rect 171 205 187 235
rect 225 205 241 235
<< pdiffcontact >>
rect 9 623 26 671
rect 40 623 56 671
rect 67 623 83 671
rect 114 623 130 671
rect 141 623 157 671
rect 171 623 187 671
rect 198 623 214 671
rect 225 623 241 671
rect 40 505 56 553
rect 67 505 83 553
rect 114 505 130 553
rect 141 505 157 553
rect 228 505 244 553
rect 255 505 271 553
<< psubstratetap >>
rect 114 175 130 192
rect 6 79 22 96
rect 34 79 50 96
rect 62 79 78 96
rect 90 79 106 96
rect 118 79 134 96
rect 146 79 162 96
rect 174 79 190 96
rect 202 79 218 96
rect 230 79 246 96
rect 258 79 274 96
<< nsubstratetap >>
rect 6 727 22 743
rect 34 727 50 743
rect 62 727 78 743
rect 90 727 106 743
rect 118 727 134 743
rect 146 727 162 743
rect 174 727 190 743
rect 202 727 218 743
rect 230 727 246 743
rect 258 727 274 743
<< metal1 >>
rect 0 782 288 792
rect 0 759 174 769
rect 252 759 288 769
rect 0 743 288 746
rect 0 727 6 743
rect 22 727 34 743
rect 50 727 62 743
rect 78 727 90 743
rect 106 727 118 743
rect 134 727 146 743
rect 162 727 174 743
rect 190 727 202 743
rect 218 727 230 743
rect 246 727 258 743
rect 274 727 288 743
rect 0 721 288 727
rect 9 671 26 721
rect 67 671 83 721
rect 93 701 211 711
rect 15 573 26 623
rect 43 613 53 623
rect 93 613 103 701
rect 120 681 184 691
rect 120 671 130 681
rect 174 671 184 681
rect 201 671 211 701
rect 43 603 103 613
rect 144 593 154 623
rect 174 613 184 623
rect 228 613 238 623
rect 174 603 238 613
rect 144 583 251 593
rect 15 563 238 573
rect 40 553 50 563
rect 145 553 157 563
rect 109 523 114 539
rect 228 553 238 563
rect 73 495 83 505
rect 73 485 180 495
rect 261 385 271 505
rect 120 365 127 379
rect 261 375 288 385
rect 261 358 271 375
rect 73 345 180 355
rect 73 335 83 345
rect 109 319 114 335
rect 46 295 56 305
rect 147 295 157 305
rect 228 295 238 328
rect 46 285 271 295
rect 13 265 235 275
rect 13 235 23 265
rect 70 245 150 255
rect 70 235 80 245
rect 114 192 130 205
rect 140 195 150 245
rect 174 235 184 265
rect 228 195 238 205
rect 140 185 238 195
rect 114 101 130 175
rect 261 101 271 285
rect 0 96 288 101
rect 0 79 6 96
rect 22 79 34 96
rect 50 79 62 96
rect 78 79 90 96
rect 106 79 118 96
rect 134 79 146 96
rect 162 79 174 96
rect 190 79 202 96
rect 218 79 230 96
rect 246 79 258 96
rect 274 79 288 96
rect 0 76 288 79
rect 0 53 288 63
rect 0 30 106 40
rect 120 30 288 40
rect 0 7 288 17
<< m2contact >>
rect 174 757 188 771
rect 238 758 252 772
rect 237 683 251 697
rect 70 367 85 381
rect 106 365 120 379
rect 174 367 188 381
rect 24 345 38 359
rect 106 28 120 42
<< metal2 >>
rect 24 359 36 799
rect 72 381 84 799
rect 175 743 187 757
rect 174 727 187 743
rect 175 381 187 727
rect 239 697 251 758
rect 24 0 36 345
rect 72 0 84 367
rect 107 42 119 365
<< labels >>
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 759 0 769 3 SDI
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 288 721 288 746 1 Vdd!
rlabel metal1 288 759 288 769 7 Q
rlabel metal1 288 782 288 792 7 ScanReturn
rlabel metal2 24 799 36 799 5 D
rlabel metal1 0 76 0 101 3 GND!
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 288 53 288 63 7 Clock
rlabel metal1 288 30 288 40 7 Test
rlabel metal1 288 7 288 17 8 nReset
rlabel metal1 288 76 288 101 7 GND!
rlabel metal2 24 0 36 0 1 D
rlabel metal1 288 375 288 385 7 M
rlabel metal2 72 0 84 0 1 Load
rlabel metal2 72 799 84 799 5 Load
<< end >>
