magic
tech c035u
timestamp 1384452322
<< nwell >>
rect 0 246 1441 323
rect 2 220 1441 246
rect 3 139 1441 220
<< polysilicon >>
rect 87 305 94 313
rect 579 305 586 313
rect 1065 305 1072 313
rect 33 206 40 214
rect 141 289 148 297
rect 168 289 175 297
rect 195 289 202 297
rect 249 293 256 301
rect 276 293 283 301
rect 303 293 310 301
rect 330 293 337 301
rect 357 293 364 301
rect 384 293 391 301
rect 411 293 418 301
rect 438 293 445 301
rect 525 206 532 214
rect 633 289 640 297
rect 660 289 667 297
rect 687 289 694 297
rect 741 293 748 301
rect 768 293 775 301
rect 795 293 802 301
rect 822 293 829 301
rect 849 293 856 301
rect 876 293 883 301
rect 903 293 910 301
rect 930 293 937 301
rect 1011 206 1018 214
rect 1119 289 1126 297
rect 1146 289 1153 297
rect 1173 289 1180 297
rect 1227 293 1234 301
rect 1254 293 1261 301
rect 1281 293 1288 301
rect 1308 293 1315 301
rect 1335 293 1342 301
rect 1362 293 1369 301
rect 1389 293 1396 301
rect 1416 293 1423 301
rect 33 134 40 148
rect 87 134 94 148
rect 141 134 148 148
rect 38 118 40 134
rect 92 118 94 134
rect 146 129 148 134
rect 168 129 175 148
rect 195 129 202 148
rect 249 134 256 148
rect 146 122 202 129
rect 146 118 148 122
rect 33 108 40 118
rect 87 108 94 118
rect 141 108 148 118
rect 168 108 175 122
rect 254 129 256 134
rect 276 129 283 148
rect 303 129 310 148
rect 330 129 337 148
rect 357 129 364 148
rect 384 129 391 148
rect 411 129 418 148
rect 438 131 445 148
rect 525 134 532 148
rect 579 134 586 148
rect 633 134 640 148
rect 436 129 445 131
rect 254 122 445 129
rect 254 118 256 122
rect 249 108 256 118
rect 276 108 283 122
rect 303 108 310 122
rect 330 108 337 122
rect 357 108 364 122
rect 384 108 391 122
rect 411 108 418 122
rect 438 108 445 122
rect 530 118 532 134
rect 584 118 586 134
rect 638 129 640 134
rect 660 129 667 148
rect 687 129 694 148
rect 741 134 748 148
rect 638 122 694 129
rect 638 118 640 122
rect 525 108 532 118
rect 579 108 586 118
rect 633 108 640 118
rect 660 108 667 122
rect 746 129 748 134
rect 768 129 775 148
rect 795 129 802 148
rect 822 129 829 148
rect 849 129 856 148
rect 876 129 883 148
rect 903 129 910 148
rect 930 131 937 148
rect 1011 134 1018 148
rect 1065 134 1072 148
rect 1119 134 1126 148
rect 928 129 937 131
rect 746 122 937 129
rect 746 118 748 122
rect 741 108 748 118
rect 768 108 775 122
rect 795 108 802 122
rect 822 108 829 122
rect 849 108 856 122
rect 876 108 883 122
rect 903 108 910 122
rect 930 108 937 122
rect 1016 118 1018 134
rect 1070 118 1072 134
rect 1124 129 1126 134
rect 1146 129 1153 148
rect 1173 129 1180 148
rect 1227 134 1234 148
rect 1124 122 1180 129
rect 1124 118 1126 122
rect 1011 108 1018 118
rect 1065 108 1072 118
rect 1119 108 1126 118
rect 1146 108 1153 122
rect 1232 129 1234 134
rect 1254 129 1261 148
rect 1281 129 1288 148
rect 1308 129 1315 148
rect 1335 129 1342 148
rect 1362 129 1369 148
rect 1389 129 1396 148
rect 1416 131 1423 148
rect 1414 129 1423 131
rect 1232 122 1423 129
rect 1232 118 1234 122
rect 1227 108 1234 118
rect 1254 108 1261 122
rect 1281 108 1288 122
rect 1308 108 1315 122
rect 1335 108 1342 122
rect 1362 108 1369 122
rect 1389 108 1396 122
rect 1416 108 1423 122
rect 33 80 40 88
rect 87 46 94 54
rect 525 80 532 88
rect 249 50 256 58
rect 276 50 283 58
rect 303 50 310 58
rect 330 50 337 58
rect 357 50 364 58
rect 384 50 391 58
rect 411 50 418 58
rect 438 50 445 58
rect 579 46 586 54
rect 1011 80 1018 88
rect 741 50 748 58
rect 768 50 775 58
rect 795 50 802 58
rect 822 50 829 58
rect 849 50 856 58
rect 876 50 883 58
rect 903 50 910 58
rect 930 50 937 58
rect 1065 46 1072 54
rect 1227 50 1234 58
rect 1254 50 1261 58
rect 1281 50 1288 58
rect 1308 50 1315 58
rect 1335 50 1342 58
rect 1362 50 1369 58
rect 1389 50 1396 58
rect 1416 50 1423 58
rect 141 27 148 35
rect 168 27 175 35
rect 633 27 640 35
rect 660 27 667 35
rect 1119 27 1126 35
rect 1146 27 1153 35
<< ndiffusion >>
rect 31 88 33 108
rect 40 88 42 108
rect 58 88 69 108
rect 85 54 87 108
rect 94 54 96 108
rect 112 54 123 108
rect 139 35 141 108
rect 148 35 150 108
rect 166 35 168 108
rect 175 35 177 108
rect 247 58 249 108
rect 256 58 258 108
rect 274 58 276 108
rect 283 58 285 108
rect 301 58 303 108
rect 310 58 312 108
rect 328 58 330 108
rect 337 58 339 108
rect 355 58 357 108
rect 364 58 366 108
rect 382 58 384 108
rect 391 58 393 108
rect 409 58 411 108
rect 418 58 420 108
rect 436 58 438 108
rect 445 58 447 108
rect 523 88 525 108
rect 532 88 534 108
rect 550 88 561 108
rect 577 54 579 108
rect 586 54 588 108
rect 604 54 615 108
rect 631 35 633 108
rect 640 35 642 108
rect 658 35 660 108
rect 667 35 669 108
rect 739 58 741 108
rect 748 58 750 108
rect 766 58 768 108
rect 775 58 777 108
rect 793 58 795 108
rect 802 58 804 108
rect 820 58 822 108
rect 829 58 831 108
rect 847 58 849 108
rect 856 58 858 108
rect 874 58 876 108
rect 883 58 885 108
rect 901 58 903 108
rect 910 58 912 108
rect 928 58 930 108
rect 937 58 939 108
rect 1009 88 1011 108
rect 1018 88 1020 108
rect 1036 88 1047 108
rect 1063 54 1065 108
rect 1072 54 1074 108
rect 1090 54 1101 108
rect 1117 35 1119 108
rect 1126 35 1128 108
rect 1144 35 1146 108
rect 1153 35 1155 108
rect 1225 58 1227 108
rect 1234 58 1236 108
rect 1252 58 1254 108
rect 1261 58 1263 108
rect 1279 58 1281 108
rect 1288 58 1290 108
rect 1306 58 1308 108
rect 1315 58 1317 108
rect 1333 58 1335 108
rect 1342 58 1344 108
rect 1360 58 1362 108
rect 1369 58 1371 108
rect 1387 58 1389 108
rect 1396 58 1398 108
rect 1414 58 1416 108
rect 1423 58 1425 108
<< pdiffusion >>
rect 31 148 33 206
rect 40 148 42 206
rect 58 148 69 206
rect 85 148 87 305
rect 94 148 96 305
rect 112 148 123 289
rect 139 148 141 289
rect 148 148 150 289
rect 166 148 168 289
rect 175 148 177 289
rect 193 148 195 289
rect 202 148 204 289
rect 220 148 231 289
rect 247 148 249 293
rect 256 148 258 293
rect 274 148 276 293
rect 283 148 285 293
rect 301 148 303 293
rect 310 148 312 293
rect 328 148 330 293
rect 337 148 339 293
rect 355 148 357 293
rect 364 148 366 293
rect 382 148 384 293
rect 391 148 393 293
rect 409 148 411 293
rect 418 148 420 293
rect 436 148 438 293
rect 445 148 447 293
rect 523 148 525 206
rect 532 148 534 206
rect 550 148 561 206
rect 577 148 579 305
rect 586 148 588 305
rect 604 148 615 289
rect 631 148 633 289
rect 640 148 642 289
rect 658 148 660 289
rect 667 148 669 289
rect 685 148 687 289
rect 694 148 696 289
rect 712 148 723 289
rect 739 148 741 293
rect 748 148 750 293
rect 766 148 768 293
rect 775 148 777 293
rect 793 148 795 293
rect 802 148 804 293
rect 820 148 822 293
rect 829 148 831 293
rect 847 148 849 293
rect 856 148 858 293
rect 874 148 876 293
rect 883 148 885 293
rect 901 148 903 293
rect 910 148 912 293
rect 928 148 930 293
rect 937 148 939 293
rect 1009 148 1011 206
rect 1018 148 1020 206
rect 1036 148 1047 206
rect 1063 148 1065 305
rect 1072 148 1074 305
rect 1090 148 1101 289
rect 1117 148 1119 289
rect 1126 148 1128 289
rect 1144 148 1146 289
rect 1153 148 1155 289
rect 1171 148 1173 289
rect 1180 148 1182 289
rect 1198 148 1209 289
rect 1225 148 1227 293
rect 1234 148 1236 293
rect 1252 148 1254 293
rect 1261 148 1263 293
rect 1279 148 1281 293
rect 1288 148 1290 293
rect 1306 148 1308 293
rect 1315 148 1317 293
rect 1333 148 1335 293
rect 1342 148 1344 293
rect 1360 148 1362 293
rect 1369 148 1371 293
rect 1387 148 1389 293
rect 1396 148 1398 293
rect 1414 148 1416 293
rect 1423 148 1425 293
<< ntransistor >>
rect 33 88 40 108
rect 87 54 94 108
rect 141 35 148 108
rect 168 35 175 108
rect 249 58 256 108
rect 276 58 283 108
rect 303 58 310 108
rect 330 58 337 108
rect 357 58 364 108
rect 384 58 391 108
rect 411 58 418 108
rect 438 58 445 108
rect 525 88 532 108
rect 579 54 586 108
rect 633 35 640 108
rect 660 35 667 108
rect 741 58 748 108
rect 768 58 775 108
rect 795 58 802 108
rect 822 58 829 108
rect 849 58 856 108
rect 876 58 883 108
rect 903 58 910 108
rect 930 58 937 108
rect 1011 88 1018 108
rect 1065 54 1072 108
rect 1119 35 1126 108
rect 1146 35 1153 108
rect 1227 58 1234 108
rect 1254 58 1261 108
rect 1281 58 1288 108
rect 1308 58 1315 108
rect 1335 58 1342 108
rect 1362 58 1369 108
rect 1389 58 1396 108
rect 1416 58 1423 108
<< ptransistor >>
rect 33 148 40 206
rect 87 148 94 305
rect 141 148 148 289
rect 168 148 175 289
rect 195 148 202 289
rect 249 148 256 293
rect 276 148 283 293
rect 303 148 310 293
rect 330 148 337 293
rect 357 148 364 293
rect 384 148 391 293
rect 411 148 418 293
rect 438 148 445 293
rect 525 148 532 206
rect 579 148 586 305
rect 633 148 640 289
rect 660 148 667 289
rect 687 148 694 289
rect 741 148 748 293
rect 768 148 775 293
rect 795 148 802 293
rect 822 148 829 293
rect 849 148 856 293
rect 876 148 883 293
rect 903 148 910 293
rect 930 148 937 293
rect 1011 148 1018 206
rect 1065 148 1072 305
rect 1119 148 1126 289
rect 1146 148 1153 289
rect 1173 148 1180 289
rect 1227 148 1234 293
rect 1254 148 1261 293
rect 1281 148 1288 293
rect 1308 148 1315 293
rect 1335 148 1342 293
rect 1362 148 1369 293
rect 1389 148 1396 293
rect 1416 148 1423 293
<< polycontact >>
rect 22 118 38 134
rect 76 118 92 134
rect 130 118 146 134
rect 238 118 254 134
rect 514 118 530 134
rect 568 118 584 134
rect 622 118 638 134
rect 730 118 746 134
rect 1000 118 1016 134
rect 1054 118 1070 134
rect 1108 118 1124 134
rect 1216 118 1232 134
<< ndiffcontact >>
rect 15 88 31 108
rect 42 88 58 108
rect 69 54 85 108
rect 96 54 112 108
rect 123 35 139 108
rect 150 35 166 108
rect 177 35 193 108
rect 231 58 247 108
rect 258 58 274 108
rect 285 58 301 108
rect 312 58 328 108
rect 339 58 355 108
rect 366 58 382 108
rect 393 58 409 108
rect 420 58 436 108
rect 447 58 463 108
rect 507 88 523 108
rect 534 88 550 108
rect 561 54 577 108
rect 588 54 604 108
rect 615 35 631 108
rect 642 35 658 108
rect 669 35 685 108
rect 723 58 739 108
rect 750 58 766 108
rect 777 58 793 108
rect 804 58 820 108
rect 831 58 847 108
rect 858 58 874 108
rect 885 58 901 108
rect 912 58 928 108
rect 939 58 955 108
rect 993 88 1009 108
rect 1020 88 1036 108
rect 1047 54 1063 108
rect 1074 54 1090 108
rect 1101 35 1117 108
rect 1128 35 1144 108
rect 1155 35 1171 108
rect 1209 58 1225 108
rect 1236 58 1252 108
rect 1263 58 1279 108
rect 1290 58 1306 108
rect 1317 58 1333 108
rect 1344 58 1360 108
rect 1371 58 1387 108
rect 1398 58 1414 108
rect 1425 58 1441 108
<< pdiffcontact >>
rect 15 148 31 206
rect 42 148 58 206
rect 69 148 85 305
rect 96 148 112 305
rect 123 148 139 289
rect 150 148 166 289
rect 177 148 193 289
rect 204 148 220 289
rect 231 148 247 293
rect 258 148 274 293
rect 285 148 301 293
rect 312 148 328 293
rect 339 148 355 293
rect 366 148 382 293
rect 393 148 409 293
rect 420 148 436 293
rect 447 148 463 293
rect 507 148 523 206
rect 534 148 550 206
rect 561 148 577 305
rect 588 148 604 305
rect 615 148 631 289
rect 642 148 658 289
rect 669 148 685 289
rect 696 148 712 289
rect 723 148 739 293
rect 750 148 766 293
rect 777 148 793 293
rect 804 148 820 293
rect 831 148 847 293
rect 858 148 874 293
rect 885 148 901 293
rect 912 148 928 293
rect 939 148 955 293
rect 993 148 1009 206
rect 1020 148 1036 206
rect 1047 148 1063 305
rect 1074 148 1090 305
rect 1101 148 1117 289
rect 1128 148 1144 289
rect 1155 148 1171 289
rect 1182 148 1198 289
rect 1209 148 1225 293
rect 1236 148 1252 293
rect 1263 148 1279 293
rect 1290 148 1306 293
rect 1317 148 1333 293
rect 1344 148 1360 293
rect 1371 148 1387 293
rect 1398 148 1414 293
rect 1425 148 1441 293
<< metal1 >>
rect -104 375 1489 385
rect -104 351 1489 361
rect -149 315 1489 340
rect 15 206 31 315
rect 69 305 85 315
rect 123 289 139 315
rect 177 289 193 315
rect 231 293 247 315
rect 285 293 301 315
rect 339 293 355 315
rect 393 293 409 315
rect 447 293 463 315
rect 507 206 523 315
rect 561 305 577 315
rect -81 119 22 129
rect 48 131 58 148
rect 48 121 76 131
rect 48 108 58 121
rect 102 131 112 148
rect 102 121 130 131
rect 102 108 112 121
rect 156 131 166 148
rect 210 131 220 148
rect 156 121 238 131
rect 156 108 166 121
rect 264 131 274 148
rect 318 131 328 148
rect 372 131 382 148
rect 426 131 436 148
rect 615 289 631 315
rect 669 289 685 315
rect 723 293 739 315
rect 777 293 793 315
rect 831 293 847 315
rect 885 293 901 315
rect 939 293 955 315
rect 993 206 1009 315
rect 1047 305 1063 315
rect 264 121 446 131
rect 264 108 274 121
rect 318 108 328 121
rect 372 108 382 121
rect 426 108 436 121
rect 476 129 486 145
rect 476 119 514 129
rect 540 131 550 148
rect 540 121 568 131
rect 540 108 550 121
rect 594 131 604 148
rect 594 121 622 131
rect 594 108 604 121
rect 648 131 658 148
rect 702 131 712 148
rect 648 121 730 131
rect 648 108 658 121
rect 756 131 766 148
rect 810 131 820 148
rect 864 131 874 148
rect 918 131 928 148
rect 756 121 944 131
rect 756 108 766 121
rect 810 108 820 121
rect 864 108 874 121
rect 918 108 928 121
rect 969 129 979 172
rect 1101 289 1117 315
rect 1155 289 1171 315
rect 1209 293 1225 315
rect 1263 293 1279 315
rect 1317 293 1333 315
rect 1371 293 1387 315
rect 1425 293 1441 315
rect 969 119 1000 129
rect 1026 131 1036 148
rect 1026 121 1054 131
rect 1026 108 1036 121
rect 1080 131 1090 148
rect 1080 121 1108 131
rect 1080 108 1090 121
rect 1134 131 1144 148
rect 1188 131 1198 148
rect 1134 121 1216 131
rect 1134 108 1144 121
rect 1242 131 1252 148
rect 1296 131 1306 148
rect 1350 131 1360 148
rect 1404 131 1414 148
rect 1242 121 1452 131
rect 1242 108 1252 121
rect 1296 108 1306 121
rect 1350 108 1360 121
rect 1404 108 1414 121
rect 15 25 31 88
rect 69 25 85 54
rect 123 25 139 35
rect 177 25 193 35
rect 231 25 247 58
rect 285 25 301 58
rect 339 25 355 58
rect 393 25 409 58
rect 447 25 463 58
rect 507 25 523 88
rect 561 25 577 54
rect 615 25 631 35
rect 669 25 685 35
rect 723 25 739 58
rect 777 25 793 58
rect 831 25 847 58
rect 885 25 901 58
rect 939 25 955 58
rect 993 25 1009 88
rect 1047 25 1063 54
rect 1101 25 1117 35
rect 1155 25 1171 35
rect 1209 25 1225 58
rect 1263 25 1279 58
rect 1317 25 1333 58
rect 1371 25 1387 58
rect 1425 25 1441 58
rect 15 0 1489 25
rect 1465 -24 1489 -14
rect 982 -44 1489 -34
rect 481 -64 1489 -54
<< m2contact >>
rect -118 374 -104 388
rect -118 350 -104 364
rect -163 315 -149 340
rect -95 119 -81 133
rect 474 145 488 159
rect 965 172 979 186
rect 446 119 460 133
rect 944 119 958 133
rect 1452 119 1466 133
rect 1451 -24 1465 -10
rect 968 -44 982 -30
rect 467 -66 481 -52
<< metal2 >>
rect -338 340 -138 422
rect -116 388 -104 422
rect -338 315 -163 340
rect -149 315 -138 340
rect -338 -78 -138 315
rect -117 -78 -105 350
rect -94 133 -82 422
rect -72 158 -60 422
rect -50 186 -38 422
rect -50 174 965 186
rect -72 146 474 158
rect 460 119 480 131
rect 958 120 980 132
rect 468 -52 480 119
rect 968 -30 980 120
rect 1452 -10 1464 119
<< end >>
