magic
tech c035u
timestamp 1385494507
<< nwell >>
rect 0 406 528 750
<< polysilicon >>
rect 44 715 51 723
rect 74 715 81 723
rect 186 715 193 723
rect 276 715 283 723
rect 331 715 338 723
rect 495 715 502 723
rect 44 130 51 667
rect 74 657 81 667
rect 74 611 81 641
rect 186 637 193 667
rect 131 611 138 619
rect 186 611 193 621
rect 276 611 283 667
rect 331 657 338 667
rect 74 533 81 563
rect 74 454 81 485
rect 74 366 81 406
rect 74 286 81 336
rect 74 226 81 256
rect 74 166 81 196
rect 74 130 81 150
rect 131 130 138 563
rect 186 533 193 563
rect 276 533 283 563
rect 186 454 193 485
rect 241 454 248 462
rect 276 437 283 485
rect 186 366 193 406
rect 241 346 248 406
rect 186 286 193 336
rect 276 339 283 421
rect 241 308 248 316
rect 276 286 283 323
rect 186 226 193 256
rect 276 226 283 256
rect 186 166 193 196
rect 186 130 193 150
rect 276 130 283 196
rect 331 176 338 641
rect 367 611 374 621
rect 394 611 401 683
rect 451 611 458 621
rect 367 553 374 563
rect 367 539 381 553
rect 394 539 401 563
rect 451 539 458 563
rect 363 500 370 508
rect 424 500 431 508
rect 451 500 458 508
rect 495 484 502 667
rect 363 422 370 452
rect 363 376 370 406
rect 424 399 431 452
rect 451 442 458 452
rect 363 329 370 360
rect 424 329 431 383
rect 451 375 458 426
rect 451 329 458 359
rect 495 352 502 468
rect 363 291 370 299
rect 424 291 431 299
rect 451 291 458 299
rect 367 236 374 260
rect 396 236 403 260
rect 451 236 458 246
rect 367 196 374 206
rect 331 130 338 160
rect 396 153 403 206
rect 451 196 458 206
rect 44 92 51 100
rect 74 92 81 100
rect 131 92 138 100
rect 186 92 193 100
rect 276 92 283 100
rect 331 92 338 100
rect 396 98 403 137
rect 495 130 502 336
rect 495 92 502 100
<< ndiffusion >>
rect 72 336 74 366
rect 81 336 83 366
rect 72 256 74 286
rect 81 256 83 286
rect 72 196 74 226
rect 81 196 83 226
rect 184 336 186 366
rect 193 336 195 366
rect 239 316 241 346
rect 248 316 250 346
rect 184 256 186 286
rect 193 256 195 286
rect 274 256 276 286
rect 283 256 285 286
rect 184 196 186 226
rect 193 196 195 226
rect 274 196 276 226
rect 283 196 285 226
rect 361 299 363 329
rect 370 299 378 329
rect 422 299 424 329
rect 431 299 433 329
rect 449 299 451 329
rect 458 299 460 329
rect 365 206 367 236
rect 374 206 378 236
rect 394 206 396 236
rect 403 206 418 236
rect 434 206 451 236
rect 458 206 460 236
rect 42 100 44 130
rect 51 100 53 130
rect 69 100 74 130
rect 81 100 85 130
rect 129 100 131 130
rect 138 100 140 130
rect 184 100 186 130
rect 193 100 202 130
rect 274 100 276 130
rect 283 100 285 130
rect 329 100 331 130
rect 338 100 340 130
rect 493 100 495 130
rect 502 100 504 130
<< pdiffusion >>
rect 42 667 44 715
rect 51 667 56 715
rect 72 667 74 715
rect 81 667 85 715
rect 184 667 186 715
rect 193 667 195 715
rect 274 667 276 715
rect 283 667 285 715
rect 329 667 331 715
rect 338 667 340 715
rect 72 563 74 611
rect 81 563 85 611
rect 129 563 131 611
rect 138 563 166 611
rect 182 563 186 611
rect 193 563 202 611
rect 274 563 276 611
rect 283 563 285 611
rect 72 485 74 533
rect 81 485 85 533
rect 72 406 74 454
rect 81 406 85 454
rect 184 485 186 533
rect 193 485 195 533
rect 274 485 276 533
rect 283 485 285 533
rect 184 406 186 454
rect 193 406 195 454
rect 211 406 241 454
rect 248 406 250 454
rect 493 667 495 715
rect 502 667 504 715
rect 363 563 367 611
rect 374 563 394 611
rect 401 563 403 611
rect 447 563 451 611
rect 458 563 460 611
rect 361 452 363 500
rect 370 452 378 500
rect 394 452 424 500
rect 431 452 451 500
rect 458 452 460 500
<< pohmic >>
rect 0 65 10 75
rect 26 65 38 75
rect 54 65 66 75
rect 82 65 94 75
rect 110 65 122 75
rect 138 65 150 75
rect 166 65 178 75
rect 194 65 206 75
rect 222 65 234 75
rect 250 65 262 75
rect 278 65 290 75
rect 306 65 318 75
rect 334 65 346 75
rect 362 65 374 75
rect 390 65 402 75
rect 418 65 430 75
rect 446 65 458 75
rect 474 65 486 75
rect 502 65 528 75
<< nohmic >>
rect 0 740 13 750
rect 29 740 41 750
rect 57 740 69 750
rect 85 740 97 750
rect 113 740 125 750
rect 141 740 153 750
rect 169 740 181 750
rect 197 740 209 750
rect 225 740 237 750
rect 253 740 265 750
rect 281 740 293 750
rect 309 740 321 750
rect 337 740 349 750
rect 365 740 377 750
rect 393 740 405 750
rect 421 740 433 750
rect 449 740 461 750
rect 477 740 489 750
rect 505 740 528 750
<< ntransistor >>
rect 74 336 81 366
rect 74 256 81 286
rect 74 196 81 226
rect 186 336 193 366
rect 241 316 248 346
rect 186 256 193 286
rect 276 256 283 286
rect 186 196 193 226
rect 276 196 283 226
rect 363 299 370 329
rect 424 299 431 329
rect 451 299 458 329
rect 367 206 374 236
rect 396 206 403 236
rect 451 206 458 236
rect 44 100 51 130
rect 74 100 81 130
rect 131 100 138 130
rect 186 100 193 130
rect 276 100 283 130
rect 331 100 338 130
rect 495 100 502 130
<< ptransistor >>
rect 44 667 51 715
rect 74 667 81 715
rect 186 667 193 715
rect 276 667 283 715
rect 331 667 338 715
rect 74 563 81 611
rect 131 563 138 611
rect 186 563 193 611
rect 276 563 283 611
rect 74 485 81 533
rect 74 406 81 454
rect 186 485 193 533
rect 276 485 283 533
rect 186 406 193 454
rect 241 406 248 454
rect 495 667 502 715
rect 367 563 374 611
rect 394 563 401 611
rect 451 563 458 611
rect 363 452 370 500
rect 424 452 431 500
rect 451 452 458 500
<< polycontact >>
rect 390 683 406 699
rect 65 641 81 657
rect 182 621 198 637
rect 326 641 342 657
rect 65 150 81 166
rect 276 421 292 437
rect 276 323 292 339
rect 181 150 197 166
rect 363 621 379 637
rect 446 621 462 637
rect 486 468 502 484
rect 358 406 374 422
rect 446 426 462 442
rect 418 383 434 399
rect 358 360 374 376
rect 446 359 462 375
rect 486 336 502 352
rect 358 180 374 196
rect 326 160 342 176
rect 446 180 462 196
rect 390 137 406 153
<< ndiffcontact >>
rect 56 336 72 366
rect 83 336 99 366
rect 56 256 72 286
rect 83 256 99 286
rect 56 196 72 226
rect 83 196 99 226
rect 168 336 184 366
rect 195 336 211 366
rect 223 316 239 346
rect 250 316 266 346
rect 168 256 184 286
rect 195 256 211 286
rect 258 256 274 286
rect 285 256 301 286
rect 168 196 184 226
rect 195 196 211 226
rect 258 196 274 226
rect 285 196 301 226
rect 345 299 361 329
rect 378 299 394 329
rect 406 299 422 329
rect 433 299 449 329
rect 460 299 476 329
rect 347 206 365 236
rect 378 206 394 236
rect 418 206 434 236
rect 460 206 476 236
rect 26 100 42 130
rect 53 100 69 130
rect 85 100 101 130
rect 113 100 129 130
rect 140 100 156 130
rect 168 100 184 130
rect 202 100 218 130
rect 258 100 274 130
rect 285 100 301 130
rect 313 100 329 130
rect 340 100 356 130
rect 477 100 493 130
rect 504 100 520 130
<< pdiffcontact >>
rect 26 667 42 715
rect 56 667 72 715
rect 85 667 101 715
rect 168 667 184 715
rect 195 667 211 715
rect 258 667 274 715
rect 285 667 301 715
rect 313 667 329 715
rect 340 667 356 715
rect 56 563 72 611
rect 85 563 101 611
rect 113 563 129 611
rect 166 563 182 611
rect 202 563 218 611
rect 258 563 274 611
rect 285 563 301 611
rect 56 485 72 533
rect 85 485 101 533
rect 56 406 72 454
rect 85 406 101 454
rect 168 485 184 533
rect 195 485 211 533
rect 258 485 274 533
rect 285 485 301 533
rect 168 406 184 454
rect 195 406 211 454
rect 250 406 266 454
rect 477 667 493 715
rect 504 667 520 715
rect 347 563 363 611
rect 403 563 419 611
rect 431 563 447 611
rect 460 563 476 611
rect 345 452 361 500
rect 378 452 394 500
rect 460 452 476 500
<< psubstratetap >>
rect 10 65 26 81
rect 38 65 54 81
rect 66 65 82 81
rect 94 65 110 81
rect 122 65 138 81
rect 150 65 166 81
rect 178 65 194 81
rect 206 65 222 81
rect 234 65 250 81
rect 262 65 278 81
rect 290 65 306 81
rect 318 65 334 81
rect 346 65 362 81
rect 374 65 390 81
rect 402 65 418 81
rect 430 65 446 81
rect 458 65 474 81
rect 486 65 502 81
<< nsubstratetap >>
rect 13 734 29 750
rect 41 734 57 750
rect 69 734 85 750
rect 97 734 113 750
rect 125 734 141 750
rect 153 734 169 750
rect 181 734 197 750
rect 209 734 225 750
rect 237 734 253 750
rect 265 734 281 750
rect 293 734 309 750
rect 321 734 337 750
rect 349 734 365 750
rect 377 734 393 750
rect 405 734 421 750
rect 433 734 449 750
rect 461 734 477 750
rect 489 734 505 750
<< metal1 >>
rect 0 780 528 790
rect 0 760 528 770
rect 0 734 13 750
rect 29 734 41 750
rect 57 734 69 750
rect 85 734 97 750
rect 113 734 125 750
rect 141 734 153 750
rect 169 734 181 750
rect 197 734 209 750
rect 225 734 237 750
rect 253 734 265 750
rect 281 734 293 750
rect 309 734 321 750
rect 337 734 349 750
rect 365 734 377 750
rect 393 734 405 750
rect 421 734 433 750
rect 449 734 461 750
rect 477 734 489 750
rect 505 734 528 750
rect 0 725 528 734
rect 6 553 16 725
rect 59 715 69 725
rect 316 715 326 725
rect 507 715 517 725
rect 101 686 168 696
rect 211 686 258 696
rect 356 686 390 696
rect 406 686 453 696
rect 467 686 477 696
rect 29 654 39 667
rect 29 644 65 654
rect 91 647 278 657
rect 91 611 101 647
rect 116 624 182 634
rect 116 611 126 624
rect 208 611 218 647
rect 268 631 278 647
rect 288 654 298 667
rect 288 644 326 654
rect 445 647 486 657
rect 268 621 363 631
rect 406 621 446 631
rect 288 611 298 621
rect 406 611 416 621
rect 476 601 486 647
rect 59 553 69 563
rect 116 553 126 563
rect 169 553 179 563
rect 260 553 270 563
rect 347 553 357 563
rect 6 543 357 553
rect 59 533 69 543
rect 260 533 270 543
rect 101 504 168 514
rect 211 504 238 514
rect 59 475 69 485
rect 228 475 238 504
rect 347 520 357 543
rect 431 520 441 563
rect 301 504 333 514
rect 347 510 441 520
rect 323 481 333 504
rect 381 500 391 510
rect 59 465 208 475
rect 228 465 312 475
rect 323 471 345 481
rect 59 454 69 465
rect 198 454 208 465
rect 101 425 168 435
rect 148 396 158 425
rect 266 425 276 435
rect 302 416 312 465
rect 476 471 486 481
rect 348 442 358 452
rect 348 432 446 442
rect 302 406 358 416
rect 148 386 418 396
rect 198 366 208 386
rect 99 342 168 352
rect 302 366 358 376
rect 59 326 69 336
rect 59 316 223 326
rect 266 326 276 336
rect 59 286 69 316
rect 302 306 312 366
rect 384 359 446 369
rect 384 329 394 359
rect 409 339 486 349
rect 409 329 419 339
rect 463 329 473 339
rect 123 296 312 306
rect 323 309 345 319
rect 123 276 133 296
rect 99 266 168 276
rect 323 276 333 309
rect 436 289 446 299
rect 301 266 333 276
rect 347 279 446 289
rect 59 246 69 256
rect 198 246 208 256
rect 261 246 271 256
rect 347 246 357 279
rect 6 236 357 246
rect 421 236 431 279
rect 6 90 16 236
rect 59 226 69 236
rect 99 206 168 216
rect 211 206 258 216
rect 301 206 321 216
rect 311 196 321 206
rect 384 196 394 206
rect 311 186 358 196
rect 91 176 298 186
rect 384 186 446 196
rect 29 153 65 163
rect 29 130 39 153
rect 91 130 101 176
rect 143 153 181 163
rect 143 130 153 153
rect 208 130 218 176
rect 288 166 326 176
rect 288 130 298 166
rect 316 140 390 150
rect 316 130 326 140
rect 476 164 486 216
rect 442 154 486 164
rect 356 110 453 120
rect 467 110 477 120
rect 56 90 66 100
rect 116 90 126 100
rect 171 90 181 100
rect 261 90 271 100
rect 507 90 517 100
rect 0 81 528 90
rect 0 65 10 81
rect 26 65 38 81
rect 54 65 66 81
rect 82 65 94 81
rect 110 65 122 81
rect 138 65 150 81
rect 166 65 178 81
rect 194 65 206 81
rect 222 65 234 81
rect 250 65 262 81
rect 278 65 290 81
rect 306 65 318 81
rect 334 65 346 81
rect 362 65 374 81
rect 390 65 402 81
rect 418 65 430 81
rect 446 65 458 81
rect 474 65 486 81
rect 502 65 528 81
rect 0 45 528 55
rect 0 25 528 35
rect 0 5 528 15
<< m2contact >>
rect 453 683 467 698
rect 431 647 445 661
rect 367 539 381 553
rect 392 539 406 553
rect 451 539 465 553
rect 43 382 57 396
rect 128 362 142 376
rect 237 362 251 376
rect 367 246 381 260
rect 392 246 406 260
rect 451 246 465 260
rect 428 152 442 166
rect 453 108 467 122
<< metal2 >>
rect 48 396 60 795
rect 57 382 60 396
rect 48 0 60 382
rect 120 376 132 795
rect 240 376 252 795
rect 432 720 444 795
rect 430 708 444 720
rect 430 661 442 708
rect 456 698 468 795
rect 467 695 468 698
rect 467 683 514 695
rect 430 659 431 661
rect 120 362 128 376
rect 251 362 252 376
rect 120 0 132 362
rect 240 0 252 362
rect 343 647 431 659
rect 343 166 355 647
rect 368 260 380 539
rect 393 260 405 539
rect 452 260 464 539
rect 343 154 428 166
rect 429 98 441 152
rect 467 120 468 122
rect 502 120 514 683
rect 467 108 514 120
rect 429 86 444 98
rect 432 0 444 86
rect 456 0 468 108
<< labels >>
rlabel metal1 0 780 0 790 3 ScanReturn
rlabel metal1 0 760 0 770 3 Q
rlabel metal1 0 725 0 750 3 Vdd!
rlabel metal1 528 780 528 790 7 ScanReturn
rlabel metal1 528 760 528 770 7 Q
rlabel metal1 528 725 528 750 7 Vdd!
rlabel metal1 0 65 0 90 3 GND!
rlabel metal1 0 45 0 55 3 Clock
rlabel metal1 0 25 0 35 3 Test
rlabel metal1 0 5 0 15 3 Reset
rlabel metal1 528 65 528 90 7 GND!
rlabel metal1 528 45 528 55 7 Clock
rlabel metal1 528 25 528 35 7 Test
rlabel metal1 528 5 528 15 7 Reset
rlabel metal2 456 0 468 0 1 Cout
rlabel metal2 432 0 444 0 1 S
rlabel metal2 240 0 252 0 1 Cin
rlabel metal2 120 0 132 0 1 B
rlabel metal2 48 0 60 0 1 A
rlabel metal2 48 795 60 795 5 A
rlabel metal2 120 795 132 795 5 B
rlabel metal2 240 795 252 795 5 Cin
rlabel metal2 432 795 444 795 5 S
rlabel metal2 456 795 468 795 5 Cout
<< end >>
