magic
tech c035u
timestamp 1384600137
<< nwell >>
rect 18 473 348 793
rect 14 415 349 473
<< polysilicon >>
rect 37 669 44 802
rect 68 761 75 802
rect 99 761 106 802
rect 37 203 44 621
rect 68 527 75 713
rect 99 670 106 713
rect 135 670 142 802
rect 176 670 183 802
rect 212 787 219 802
rect 212 757 219 771
rect 250 757 257 802
rect 212 670 219 709
rect 99 527 106 622
rect 135 527 142 622
rect 176 605 183 622
rect 176 527 183 589
rect 212 527 219 622
rect 250 579 257 709
rect 282 607 289 802
rect 323 787 330 802
rect 323 670 330 771
rect 68 313 75 479
rect 99 373 106 479
rect 135 469 142 479
rect 135 373 142 453
rect 99 313 106 325
rect 37 55 44 155
rect 68 143 75 265
rect 99 203 106 265
rect 135 203 142 325
rect 176 313 183 479
rect 212 469 219 479
rect 212 313 219 453
rect 176 171 183 265
rect 212 229 219 265
rect 212 203 219 213
rect 250 203 257 563
rect 282 527 289 591
rect 282 347 289 479
rect 323 373 330 622
rect 282 313 289 331
rect 68 55 75 95
rect 99 55 106 155
rect 135 79 142 155
rect 176 143 183 155
rect 212 143 219 155
rect 250 143 257 155
rect 135 55 142 63
rect 176 53 183 95
rect 212 53 219 95
rect 250 55 257 95
rect 282 55 289 265
rect 323 203 330 325
rect 323 55 330 155
<< ndiffusion >>
rect 97 325 99 373
rect 106 325 135 373
rect 142 325 149 373
rect 66 265 68 313
rect 75 265 99 313
rect 106 265 114 313
rect 35 155 37 203
rect 44 155 46 203
rect 173 265 176 313
rect 183 265 212 313
rect 219 265 224 313
rect 97 155 99 203
rect 106 155 135 203
rect 142 155 146 203
rect 317 325 323 373
rect 330 325 340 373
rect 280 265 282 313
rect 289 265 295 313
rect 209 155 212 203
rect 219 155 250 203
rect 257 155 261 203
rect 66 95 68 143
rect 75 95 78 143
rect 171 95 176 143
rect 183 95 212 143
rect 219 95 223 143
<< pdiffusion >>
rect 65 713 68 761
rect 75 713 78 761
rect 94 713 99 761
rect 106 713 108 761
rect 34 621 37 669
rect 44 621 46 669
rect 209 709 212 757
rect 219 709 229 757
rect 245 709 250 757
rect 257 709 260 757
rect 96 622 99 670
rect 106 622 110 670
rect 126 622 135 670
rect 142 622 155 670
rect 173 622 176 670
rect 183 622 193 670
rect 209 622 212 670
rect 219 622 221 670
rect 320 622 323 670
rect 330 622 332 670
rect 65 479 68 527
rect 75 479 80 527
rect 96 479 99 527
rect 106 479 109 527
rect 125 479 135 527
rect 142 479 155 527
rect 173 479 176 527
rect 183 479 185 527
rect 201 479 212 527
rect 219 479 222 527
rect 279 479 282 527
rect 289 479 291 527
<< ntransistor >>
rect 99 325 106 373
rect 135 325 142 373
rect 68 265 75 313
rect 99 265 106 313
rect 37 155 44 203
rect 176 265 183 313
rect 212 265 219 313
rect 99 155 106 203
rect 135 155 142 203
rect 323 325 330 373
rect 282 265 289 313
rect 212 155 219 203
rect 250 155 257 203
rect 68 95 75 143
rect 176 95 183 143
rect 212 95 219 143
<< ptransistor >>
rect 68 713 75 761
rect 99 713 106 761
rect 37 621 44 669
rect 212 709 219 757
rect 250 709 257 757
rect 99 622 106 670
rect 135 622 142 670
rect 176 622 183 670
rect 212 622 219 670
rect 323 622 330 670
rect 68 479 75 527
rect 99 479 106 527
rect 135 479 142 527
rect 176 479 183 527
rect 212 479 219 527
rect 282 479 289 527
<< polycontact >>
rect 203 771 219 787
rect 167 589 183 605
rect 314 771 330 787
rect 273 591 289 607
rect 245 563 261 579
rect 130 453 146 469
rect 212 453 228 469
rect 212 213 228 229
rect 273 331 289 347
rect 167 155 183 171
rect 250 95 266 143
rect 135 63 151 79
rect 314 155 330 203
<< ndiffcontact >>
rect 81 325 97 373
rect 149 325 165 373
rect 50 265 66 313
rect 114 265 130 313
rect 19 155 35 203
rect 46 155 62 203
rect 157 265 173 313
rect 224 265 240 313
rect 81 155 97 203
rect 146 155 162 203
rect 301 325 317 373
rect 340 325 356 373
rect 264 265 280 313
rect 295 265 311 313
rect 193 155 209 203
rect 261 155 277 203
rect 50 95 66 143
rect 78 95 94 143
rect 155 95 171 143
rect 223 95 239 143
<< pdiffcontact >>
rect 49 713 65 761
rect 78 713 94 761
rect 108 713 124 761
rect 18 621 34 669
rect 46 621 62 669
rect 193 709 209 757
rect 229 709 245 757
rect 260 709 276 757
rect 80 622 96 670
rect 110 622 126 670
rect 155 622 173 670
rect 193 622 209 670
rect 221 622 237 670
rect 294 622 320 670
rect 332 622 348 670
rect 49 479 65 527
rect 80 479 96 527
rect 109 479 125 527
rect 155 479 173 527
rect 185 479 201 527
rect 222 479 238 527
rect 263 479 279 527
rect 291 479 307 527
<< psubstratetap >>
rect 111 387 129 403
<< nsubstratetap >>
rect 112 424 130 440
<< metal1 >>
rect 78 771 203 787
rect 229 771 314 787
rect 78 761 94 771
rect 229 757 245 771
rect 49 699 65 713
rect 108 699 124 713
rect 193 699 209 709
rect 260 699 276 709
rect 18 680 320 699
rect 18 669 34 680
rect 80 670 96 680
rect 155 670 173 680
rect 221 670 237 680
rect 18 553 34 621
rect 294 670 320 680
rect 46 605 62 621
rect 111 605 123 622
rect 193 607 209 622
rect 46 589 167 605
rect 193 591 273 607
rect 332 579 348 622
rect 109 563 245 579
rect 261 563 348 579
rect 18 537 96 553
rect 18 443 34 537
rect 80 527 96 537
rect 109 527 125 563
rect 155 537 348 553
rect 155 527 173 537
rect 222 527 238 537
rect 263 527 279 537
rect 49 469 65 479
rect 185 469 201 479
rect 291 469 307 479
rect 49 453 130 469
rect 146 453 201 469
rect 228 453 307 469
rect 332 443 348 537
rect 0 440 363 443
rect 0 424 112 440
rect 130 424 363 440
rect 0 418 363 424
rect 0 403 363 408
rect 0 387 111 403
rect 129 387 363 403
rect 0 383 363 387
rect 19 229 35 383
rect 81 373 97 383
rect 114 313 130 383
rect 165 357 301 373
rect 224 331 273 347
rect 224 313 240 331
rect 130 265 157 313
rect 50 255 66 265
rect 264 255 280 265
rect 50 239 280 255
rect 295 229 311 265
rect 19 213 193 229
rect 228 213 311 229
rect 19 203 35 213
rect 62 155 81 203
rect 177 187 193 213
rect 162 155 167 171
rect 277 155 314 203
rect 19 143 35 155
rect 340 143 356 325
rect 19 95 50 143
rect 94 95 155 143
rect 266 95 356 143
rect 223 79 239 95
rect 151 63 239 79
<< labels >>
rlabel metal1 0 383 0 408 3 GND!
rlabel metal1 0 418 0 443 3 Vdd!
rlabel polysilicon 37 802 44 802 5 D
rlabel polysilicon 68 802 75 802 5 Clk
rlabel polysilicon 99 802 106 802 5 nRst
rlabel polysilicon 135 802 142 802 5 Z
rlabel polysilicon 176 802 183 802 5 W
rlabel polysilicon 212 802 219 802 5 Y
rlabel polysilicon 250 802 257 802 5 nQ
rlabel polysilicon 282 802 289 802 5 X
rlabel polysilicon 323 802 330 802 5 Q
rlabel metal1 363 383 363 408 7 GND!
rlabel metal1 363 418 363 443 7 Vdd!
<< end >>
