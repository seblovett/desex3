magic
tech c035u
timestamp 1384428762
<< nwell >>
rect 0 246 463 323
rect 2 220 463 246
rect 3 139 463 220
<< polysilicon >>
rect 87 305 94 313
rect 33 206 40 214
rect 141 289 148 297
rect 168 289 175 297
rect 195 289 202 297
rect 249 293 256 301
rect 276 293 283 301
rect 303 293 310 301
rect 330 293 337 301
rect 357 293 364 301
rect 384 293 391 301
rect 411 293 418 301
rect 438 293 445 301
rect 33 134 40 148
rect 87 134 94 148
rect 141 134 148 148
rect 38 118 40 134
rect 92 118 94 134
rect 146 129 148 134
rect 168 129 175 148
rect 195 129 202 148
rect 249 134 256 148
rect 146 122 202 129
rect 146 118 148 122
rect 33 108 40 118
rect 87 108 94 118
rect 141 108 148 118
rect 168 108 175 122
rect 254 129 256 134
rect 276 129 283 148
rect 303 129 310 148
rect 330 129 337 148
rect 357 129 364 148
rect 384 129 391 148
rect 411 129 418 148
rect 438 131 445 148
rect 436 129 445 131
rect 254 122 445 129
rect 254 118 256 122
rect 249 108 256 118
rect 276 108 283 122
rect 303 108 310 122
rect 330 108 337 122
rect 357 108 364 122
rect 384 108 391 122
rect 411 108 418 122
rect 438 108 445 122
rect 33 80 40 88
rect 87 46 94 54
rect 249 50 256 58
rect 276 50 283 58
rect 303 50 310 58
rect 330 50 337 58
rect 357 50 364 58
rect 384 50 391 58
rect 411 50 418 58
rect 438 50 445 58
rect 141 27 148 35
rect 168 27 175 35
<< ndiffusion >>
rect 31 88 33 108
rect 40 88 42 108
rect 58 88 69 108
rect 85 54 87 108
rect 94 54 96 108
rect 112 54 123 108
rect 139 35 141 108
rect 148 35 150 108
rect 166 35 168 108
rect 175 35 177 108
rect 247 58 249 108
rect 256 58 258 108
rect 274 58 276 108
rect 283 58 285 108
rect 301 58 303 108
rect 310 58 312 108
rect 328 58 330 108
rect 337 58 339 108
rect 355 58 357 108
rect 364 58 366 108
rect 382 58 384 108
rect 391 58 393 108
rect 409 58 411 108
rect 418 58 420 108
rect 436 58 438 108
rect 445 58 447 108
<< pdiffusion >>
rect 31 148 33 206
rect 40 148 42 206
rect 58 148 69 206
rect 85 148 87 305
rect 94 148 96 305
rect 112 148 123 289
rect 139 148 141 289
rect 148 148 150 289
rect 166 148 168 289
rect 175 148 177 289
rect 193 148 195 289
rect 202 148 204 289
rect 220 148 231 289
rect 247 148 249 293
rect 256 148 258 293
rect 274 148 276 293
rect 283 148 285 293
rect 301 148 303 293
rect 310 148 312 293
rect 328 148 330 293
rect 337 148 339 293
rect 355 148 357 293
rect 364 148 366 293
rect 382 148 384 293
rect 391 148 393 293
rect 409 148 411 293
rect 418 148 420 293
rect 436 148 438 293
rect 445 148 447 293
<< ntransistor >>
rect 33 88 40 108
rect 87 54 94 108
rect 141 35 148 108
rect 168 35 175 108
rect 249 58 256 108
rect 276 58 283 108
rect 303 58 310 108
rect 330 58 337 108
rect 357 58 364 108
rect 384 58 391 108
rect 411 58 418 108
rect 438 58 445 108
<< ptransistor >>
rect 33 148 40 206
rect 87 148 94 305
rect 141 148 148 289
rect 168 148 175 289
rect 195 148 202 289
rect 249 148 256 293
rect 276 148 283 293
rect 303 148 310 293
rect 330 148 337 293
rect 357 148 364 293
rect 384 148 391 293
rect 411 148 418 293
rect 438 148 445 293
<< polycontact >>
rect 22 118 38 134
rect 76 118 92 134
rect 130 118 146 134
rect 238 118 254 134
<< ndiffcontact >>
rect 15 88 31 108
rect 42 88 58 108
rect 69 54 85 108
rect 96 54 112 108
rect 123 35 139 108
rect 150 35 166 108
rect 177 35 193 108
rect 231 58 247 108
rect 258 58 274 108
rect 285 58 301 108
rect 312 58 328 108
rect 339 58 355 108
rect 366 58 382 108
rect 393 58 409 108
rect 420 58 436 108
rect 447 58 463 108
<< pdiffcontact >>
rect 15 148 31 206
rect 42 148 58 206
rect 69 148 85 305
rect 96 148 112 305
rect 123 148 139 289
rect 150 148 166 289
rect 177 148 193 289
rect 204 148 220 289
rect 231 148 247 293
rect 258 148 274 293
rect 285 148 301 293
rect 312 148 328 293
rect 339 148 355 293
rect 366 148 382 293
rect 393 148 409 293
rect 420 148 436 293
rect 447 148 463 293
<< metal1 >>
rect 1 315 464 340
rect 15 206 31 315
rect 69 305 85 315
rect 123 289 139 315
rect 177 289 193 315
rect 231 293 247 315
rect 285 293 301 315
rect 339 293 355 315
rect 393 293 409 315
rect 447 293 463 315
rect 0 119 22 129
rect 48 131 58 148
rect 48 121 76 131
rect 48 108 58 121
rect 102 131 112 148
rect 102 121 130 131
rect 102 108 112 121
rect 156 131 166 148
rect 210 131 220 148
rect 156 121 238 131
rect 156 108 166 121
rect 264 131 274 148
rect 318 131 328 148
rect 372 131 382 148
rect 426 131 436 148
rect 264 121 457 131
rect 264 108 274 121
rect 318 108 328 121
rect 372 108 382 121
rect 426 108 436 121
rect 15 25 31 88
rect 69 25 85 54
rect 123 25 139 35
rect 177 25 193 35
rect 231 25 247 58
rect 285 25 301 58
rect 339 25 355 58
rect 393 25 409 58
rect 447 25 463 58
rect 0 0 463 25
<< end >>
