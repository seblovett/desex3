magic
tech c035u
timestamp 1385926514
<< error_s >>
rect 2544 782 2548 792
rect 2736 782 2742 792
rect 2544 759 2548 769
rect 2544 402 2566 746
rect 2736 402 2760 746
rect 3872 730 3882 736
rect 2544 86 2548 101
rect 2736 96 2742 101
rect 2544 76 2550 86
rect 2736 76 2744 96
rect 3872 76 3874 92
rect 2544 53 2548 63
rect 2736 53 2742 63
rect 2544 30 2548 40
rect 2736 30 2742 40
rect 2544 7 2548 17
rect 2736 7 2742 17
use ../leftbuf/leftbuf leftbuf_0
timestamp 1385752733
transform 1 0 0 0 1 10
box 0 -10 1464 789
use ../and2/and2 and2_0
timestamp 1385636468
transform 1 0 1464 0 1 0
box 0 0 120 799
use ../nand2/nand2 nand2_0
timestamp 1385631319
transform 1 0 1584 0 1 0
box 0 0 96 799
use ../nand3/nand3 nand3_0
timestamp 1385920731
transform 1 0 1680 0 1 0
box 0 0 120 799
use ../nand4/nand4 nand4_0
timestamp 1385636690
transform 1 0 1800 0 1 0
box 0 0 144 799
use ../nor2/nor2 nor2_0
timestamp 1385632928
transform 1 0 1944 0 1 0
box 0 0 120 799
use ../nor3/nor3 nor3_0
timestamp 1385633286
transform 1 0 2064 0 1 0
box 0 0 144 799
use ../or2/or2 or2_0
timestamp 1385633707
transform 1 0 2208 0 1 0
box 0 0 144 799
use ../mux2/mux2 mux2_0
timestamp 1385634976
transform 1 0 2352 0 1 0
box 0 0 186 799
use ../smux2/smux2 smux2_0
timestamp 1385635083
transform 1 0 2544 0 1 0
box 0 0 188 799
use ../smux3/smux3 smux3_0
timestamp 1385920319
transform 1 0 2736 0 1 0
box 0 0 288 799
use ../buffer/buffer buffer_0
timestamp 1385926514
transform 1 0 3024 0 1 -1
box 0 1 120 800
use ../inv/inv inv_0
timestamp 1385924870
transform 1 0 3144 0 1 0
box 0 0 120 799
use ../trisbuf/trisbuf trisbuf_0
timestamp 1385926402
transform 1 0 3264 0 1 0
box 0 0 192 799
use ../rdtype/rdtype rdtype_0
timestamp 1385639216
transform 1 0 3456 0 1 0
box 0 0 432 799
use ../fulladder/fulladder fulladder_0
timestamp 1385909444
transform 1 0 3866 0 1 0
box 0 0 360 799
use ../halfadder/halfadder halfadder_0
timestamp 1385925245
transform 1 0 4226 0 1 0
box 0 0 312 799
use ../xor2/xor2 xor2_0
timestamp 1385920833
transform 1 0 4538 0 1 0
box 0 0 185 799
use ../tiehigh/tiehigh tiehigh_0
timestamp 1385920028
transform 1 0 4723 0 1 0
box 0 0 34 799
use ../tielow/tielow tielow_0
timestamp 1385920082
transform 1 0 4757 0 1 -1
box 0 1 34 800
use ../rowcrosser/rowcrosser rowcrosser_0
timestamp 1385919898
transform 1 0 4791 0 1 0
box 0 0 34 799
use ../rightend/rightend rightend_0
timestamp 1385751130
transform 1 0 4825 0 1 0
box 0 0 292 799
<< end >>
