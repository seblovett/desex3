magic
tech c035u
timestamp 1386362310
<< metal1 >>
rect 0 863 237 873
rect 0 815 10 863
rect 371 860 741 870
rect 0 805 46 815
rect 838 421 863 431
rect 26 76 46 86
rect 26 31 36 76
rect 26 21 117 31
rect 444 21 548 31
rect 853 31 863 421
rect 562 21 863 31
<< m2contact >>
rect 237 859 251 873
rect 357 858 371 872
rect 741 856 755 870
rect 117 21 131 35
rect 430 19 444 33
rect 548 19 562 33
<< metal2 >>
rect 190 845 202 921
rect 238 845 250 859
rect 310 845 322 921
rect 358 845 370 858
rect 478 845 490 921
rect 550 845 562 921
rect 742 870 754 921
rect 742 845 754 856
rect 70 0 82 46
rect 118 35 130 46
rect 430 33 442 46
rect 550 33 562 46
use ../inv/inv inv_3
timestamp 1386238110
transform 1 0 46 0 1 46
box 0 0 120 799
use ../inv/inv inv_4
timestamp 1386238110
transform 1 0 166 0 1 46
box 0 0 120 799
use ../inv/inv inv_0
timestamp 1386238110
transform 1 0 286 0 1 46
box 0 0 120 799
use ../inv/inv inv_1
timestamp 1386238110
transform 1 0 406 0 1 46
box 0 0 120 799
use ../inv/inv inv_2
timestamp 1386238110
transform 1 0 526 0 1 46
box 0 0 120 799
use smux2 smux2_0
timestamp 1386234984
transform 1 0 646 0 1 46
box 0 0 192 799
<< labels >>
rlabel metal2 70 0 82 0 1 nTest
rlabel metal2 190 921 202 921 1 nSDI
rlabel metal2 742 921 754 921 5 D
rlabel metal2 478 921 490 921 5 n1
rlabel metal2 550 921 562 921 5 n2
<< end >>
