magic
tech c035u
timestamp 1385634976
<< nwell >>
rect 0 402 186 746
<< polysilicon >>
rect 29 691 36 699
rect 59 691 66 699
rect 86 691 93 699
rect 113 691 120 699
rect 144 691 151 699
rect 29 612 36 643
rect 59 599 66 643
rect 29 485 36 564
rect 29 347 36 469
rect 59 347 66 583
rect 86 500 93 643
rect 92 484 93 500
rect 86 347 93 484
rect 113 488 120 643
rect 144 633 151 643
rect 147 617 151 633
rect 113 472 116 488
rect 113 347 120 472
rect 144 393 151 617
rect 146 377 151 393
rect 29 282 36 317
rect 59 278 66 317
rect 86 309 93 317
rect 113 309 120 317
rect 144 282 151 377
rect 29 243 36 252
rect 144 244 151 252
<< ndiffusion >>
rect 27 317 29 347
rect 36 317 38 347
rect 54 317 59 347
rect 66 317 86 347
rect 93 317 95 347
rect 111 317 113 347
rect 120 317 122 347
rect 27 252 29 282
rect 36 252 38 282
rect 142 252 144 282
rect 151 252 153 282
<< pdiffusion >>
rect 27 643 29 691
rect 36 643 38 691
rect 54 643 59 691
rect 66 643 68 691
rect 84 643 86 691
rect 93 643 95 691
rect 111 643 113 691
rect 120 643 123 691
rect 139 643 144 691
rect 151 643 154 691
rect 27 564 29 612
rect 36 564 38 612
<< pohmic >>
rect 0 79 6 86
rect 22 79 34 86
rect 50 79 62 86
rect 78 79 90 86
rect 106 79 118 86
rect 134 79 146 86
rect 162 79 186 86
rect 0 76 186 79
<< nohmic >>
rect 0 743 186 746
rect 0 736 8 743
rect 24 736 36 743
rect 52 736 64 743
rect 80 736 92 743
rect 108 736 121 743
rect 137 736 149 743
rect 165 736 186 743
<< ntransistor >>
rect 29 317 36 347
rect 59 317 66 347
rect 86 317 93 347
rect 113 317 120 347
rect 29 252 36 282
rect 144 252 151 282
<< ptransistor >>
rect 29 643 36 691
rect 59 643 66 691
rect 86 643 93 691
rect 113 643 120 691
rect 144 643 151 691
rect 29 564 36 612
<< polycontact >>
rect 59 583 75 599
rect 25 469 41 485
rect 76 484 92 500
rect 131 617 147 633
rect 116 472 132 488
rect 130 377 146 393
rect 59 262 75 278
<< ndiffcontact >>
rect 11 317 27 347
rect 38 317 54 347
rect 95 317 111 347
rect 122 317 138 347
rect 11 252 27 282
rect 38 252 54 282
rect 126 252 142 282
rect 153 252 169 282
<< pdiffcontact >>
rect 11 643 27 691
rect 38 643 54 691
rect 68 643 84 691
rect 95 643 111 691
rect 123 643 139 691
rect 154 643 170 691
rect 11 564 27 612
rect 38 564 54 612
<< psubstratetap >>
rect 6 79 22 95
rect 34 79 50 95
rect 62 79 78 95
rect 90 79 106 95
rect 118 79 134 95
rect 146 79 162 95
<< nsubstratetap >>
rect 8 727 24 743
rect 36 727 52 743
rect 64 727 80 743
rect 92 727 108 743
rect 121 727 137 743
rect 149 727 165 743
<< metal1 >>
rect 0 782 186 792
rect 0 759 186 769
rect 0 743 186 746
rect 0 727 8 743
rect 24 727 36 743
rect 52 727 64 743
rect 80 727 92 743
rect 108 727 121 743
rect 137 727 149 743
rect 165 727 186 743
rect 0 721 186 727
rect 11 691 27 721
rect 41 701 108 711
rect 41 691 51 701
rect 98 691 108 701
rect 123 691 139 721
rect 11 612 27 643
rect 71 629 81 643
rect 71 619 131 629
rect 54 583 59 599
rect 157 469 167 643
rect 160 455 167 469
rect 41 380 130 390
rect 41 347 51 380
rect 73 357 135 367
rect 14 307 24 317
rect 73 307 83 357
rect 125 347 135 357
rect 14 297 83 307
rect 95 282 111 317
rect 157 282 167 455
rect 54 262 59 278
rect 95 252 126 282
rect 11 101 27 252
rect 95 101 111 252
rect 0 95 186 101
rect 0 79 6 95
rect 22 79 34 95
rect 50 79 62 95
rect 78 79 90 95
rect 106 79 118 95
rect 134 79 146 95
rect 162 79 186 95
rect 0 76 186 79
rect 0 53 186 63
rect 0 30 186 40
rect 0 7 186 17
<< m2contact >>
rect 118 488 132 502
rect 41 470 55 484
rect 77 470 91 484
rect 146 455 160 469
<< metal2 >>
rect 48 484 60 799
rect 55 470 60 484
rect 48 0 60 470
rect 72 484 84 799
rect 120 502 132 799
rect 72 470 77 484
rect 72 0 84 470
rect 120 0 132 488
rect 144 469 156 799
rect 144 455 146 469
rect 144 0 156 455
<< labels >>
rlabel metal1 0 76 0 101 1 GND!
rlabel metal1 0 7 0 17 2 nReset
rlabel metal1 0 30 0 40 3 Test
rlabel metal1 0 53 0 63 3 Clock
rlabel metal1 186 76 186 101 7 GND!
rlabel metal1 186 7 186 17 8 nReset
rlabel metal1 186 30 186 40 7 Test
rlabel metal1 186 53 186 63 7 Clock
rlabel metal2 48 0 60 0 1 S
rlabel metal2 144 0 156 0 1 Y
rlabel metal2 120 0 132 0 1 I1
rlabel metal2 72 0 84 0 1 I0
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 759 0 769 3 Scan
rlabel metal1 0 782 0 792 4 ScanReturn
rlabel metal1 186 721 186 746 7 Vdd!
rlabel metal1 186 782 186 792 6 ScanReturn
rlabel metal1 186 759 186 769 7 Scan
rlabel metal2 48 799 60 799 5 S
rlabel metal2 144 799 156 799 5 Y
rlabel metal2 120 799 132 799 5 I1
rlabel metal2 72 799 84 799 5 I0
<< end >>
