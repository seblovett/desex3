magic
tech c035u
timestamp 1385631071
<< nwell >>
rect 0 408 528 752
<< polysilicon >>
rect 44 717 51 725
rect 74 717 81 725
rect 186 717 193 725
rect 276 717 283 725
rect 331 717 338 725
rect 495 717 502 725
rect 44 132 51 669
rect 74 659 81 669
rect 74 613 81 643
rect 186 639 193 669
rect 131 613 138 621
rect 186 613 193 623
rect 276 613 283 669
rect 331 659 338 669
rect 74 535 81 565
rect 74 456 81 487
rect 74 368 81 408
rect 74 288 81 338
rect 74 228 81 258
rect 74 168 81 198
rect 74 132 81 152
rect 131 132 138 565
rect 186 535 193 565
rect 276 535 283 565
rect 186 456 193 487
rect 241 456 248 464
rect 276 439 283 487
rect 186 368 193 408
rect 241 348 248 408
rect 186 288 193 338
rect 276 341 283 423
rect 241 310 248 318
rect 276 288 283 325
rect 186 228 193 258
rect 276 228 283 258
rect 186 168 193 198
rect 186 132 193 152
rect 276 132 283 198
rect 331 178 338 643
rect 367 613 374 623
rect 394 613 401 685
rect 451 613 458 623
rect 367 555 374 565
rect 367 541 381 555
rect 394 541 401 565
rect 451 541 458 565
rect 363 502 370 510
rect 424 502 431 510
rect 451 502 458 510
rect 495 486 502 669
rect 363 424 370 454
rect 363 378 370 408
rect 424 401 431 454
rect 451 444 458 454
rect 363 331 370 362
rect 424 331 431 385
rect 451 377 458 428
rect 451 331 458 361
rect 495 354 502 470
rect 363 293 370 301
rect 424 293 431 301
rect 451 293 458 301
rect 367 238 374 262
rect 396 238 403 262
rect 451 238 458 248
rect 367 198 374 208
rect 331 132 338 162
rect 396 155 403 208
rect 451 198 458 208
rect 44 94 51 102
rect 74 94 81 102
rect 131 94 138 102
rect 186 94 193 102
rect 276 94 283 102
rect 331 94 338 102
rect 396 100 403 139
rect 495 132 502 338
rect 495 94 502 102
<< ndiffusion >>
rect 72 338 74 368
rect 81 338 83 368
rect 72 258 74 288
rect 81 258 83 288
rect 72 198 74 228
rect 81 198 83 228
rect 184 338 186 368
rect 193 338 195 368
rect 239 318 241 348
rect 248 318 250 348
rect 184 258 186 288
rect 193 258 195 288
rect 274 258 276 288
rect 283 258 285 288
rect 184 198 186 228
rect 193 198 195 228
rect 274 198 276 228
rect 283 198 285 228
rect 361 301 363 331
rect 370 301 378 331
rect 422 301 424 331
rect 431 301 433 331
rect 449 301 451 331
rect 458 301 460 331
rect 365 208 367 238
rect 374 208 378 238
rect 394 208 396 238
rect 403 208 418 238
rect 434 208 451 238
rect 458 208 460 238
rect 42 102 44 132
rect 51 102 53 132
rect 69 102 74 132
rect 81 102 85 132
rect 129 102 131 132
rect 138 102 140 132
rect 184 102 186 132
rect 193 102 202 132
rect 274 102 276 132
rect 283 102 285 132
rect 329 102 331 132
rect 338 102 340 132
rect 493 102 495 132
rect 502 102 504 132
<< pdiffusion >>
rect 42 669 44 717
rect 51 669 56 717
rect 72 669 74 717
rect 81 669 85 717
rect 184 669 186 717
rect 193 669 195 717
rect 274 669 276 717
rect 283 669 285 717
rect 329 669 331 717
rect 338 669 340 717
rect 72 565 74 613
rect 81 565 85 613
rect 129 565 131 613
rect 138 565 166 613
rect 182 565 186 613
rect 193 565 202 613
rect 274 565 276 613
rect 283 565 285 613
rect 72 487 74 535
rect 81 487 85 535
rect 72 408 74 456
rect 81 408 85 456
rect 184 487 186 535
rect 193 487 195 535
rect 274 487 276 535
rect 283 487 285 535
rect 184 408 186 456
rect 193 408 195 456
rect 211 408 241 456
rect 248 408 250 456
rect 493 669 495 717
rect 502 669 504 717
rect 363 565 367 613
rect 374 565 394 613
rect 401 565 403 613
rect 447 565 451 613
rect 458 565 460 613
rect 361 454 363 502
rect 370 454 378 502
rect 394 454 424 502
rect 431 454 451 502
rect 458 454 460 502
<< pohmic >>
rect 0 67 10 77
rect 26 67 38 77
rect 54 67 66 77
rect 82 67 94 77
rect 110 67 122 77
rect 138 67 150 77
rect 166 67 178 77
rect 194 67 206 77
rect 222 67 234 77
rect 250 67 262 77
rect 278 67 290 77
rect 306 67 318 77
rect 334 67 346 77
rect 362 67 374 77
rect 390 67 402 77
rect 418 67 430 77
rect 446 67 458 77
rect 474 67 486 77
rect 502 67 528 77
<< nohmic >>
rect 0 742 13 752
rect 29 742 41 752
rect 57 742 69 752
rect 85 742 97 752
rect 113 742 125 752
rect 141 742 153 752
rect 169 742 181 752
rect 197 742 209 752
rect 225 742 237 752
rect 253 742 265 752
rect 281 742 293 752
rect 309 742 321 752
rect 337 742 349 752
rect 365 742 377 752
rect 393 742 405 752
rect 421 742 433 752
rect 449 742 461 752
rect 477 742 489 752
rect 505 742 528 752
<< ntransistor >>
rect 74 338 81 368
rect 74 258 81 288
rect 74 198 81 228
rect 186 338 193 368
rect 241 318 248 348
rect 186 258 193 288
rect 276 258 283 288
rect 186 198 193 228
rect 276 198 283 228
rect 363 301 370 331
rect 424 301 431 331
rect 451 301 458 331
rect 367 208 374 238
rect 396 208 403 238
rect 451 208 458 238
rect 44 102 51 132
rect 74 102 81 132
rect 131 102 138 132
rect 186 102 193 132
rect 276 102 283 132
rect 331 102 338 132
rect 495 102 502 132
<< ptransistor >>
rect 44 669 51 717
rect 74 669 81 717
rect 186 669 193 717
rect 276 669 283 717
rect 331 669 338 717
rect 74 565 81 613
rect 131 565 138 613
rect 186 565 193 613
rect 276 565 283 613
rect 74 487 81 535
rect 74 408 81 456
rect 186 487 193 535
rect 276 487 283 535
rect 186 408 193 456
rect 241 408 248 456
rect 495 669 502 717
rect 367 565 374 613
rect 394 565 401 613
rect 451 565 458 613
rect 363 454 370 502
rect 424 454 431 502
rect 451 454 458 502
<< polycontact >>
rect 390 685 406 701
rect 65 643 81 659
rect 182 623 198 639
rect 326 643 342 659
rect 65 152 81 168
rect 276 423 292 439
rect 276 325 292 341
rect 181 152 197 168
rect 363 623 379 639
rect 446 623 462 639
rect 486 470 502 486
rect 358 408 374 424
rect 446 428 462 444
rect 418 385 434 401
rect 358 362 374 378
rect 446 361 462 377
rect 486 338 502 354
rect 358 182 374 198
rect 326 162 342 178
rect 446 182 462 198
rect 390 139 406 155
<< ndiffcontact >>
rect 56 338 72 368
rect 83 338 99 368
rect 56 258 72 288
rect 83 258 99 288
rect 56 198 72 228
rect 83 198 99 228
rect 168 338 184 368
rect 195 338 211 368
rect 223 318 239 348
rect 250 318 266 348
rect 168 258 184 288
rect 195 258 211 288
rect 258 258 274 288
rect 285 258 301 288
rect 168 198 184 228
rect 195 198 211 228
rect 258 198 274 228
rect 285 198 301 228
rect 345 301 361 331
rect 378 301 394 331
rect 406 301 422 331
rect 433 301 449 331
rect 460 301 476 331
rect 347 208 365 238
rect 378 208 394 238
rect 418 208 434 238
rect 460 208 476 238
rect 26 102 42 132
rect 53 102 69 132
rect 85 102 101 132
rect 113 102 129 132
rect 140 102 156 132
rect 168 102 184 132
rect 202 102 218 132
rect 258 102 274 132
rect 285 102 301 132
rect 313 102 329 132
rect 340 102 356 132
rect 477 102 493 132
rect 504 102 520 132
<< pdiffcontact >>
rect 26 669 42 717
rect 56 669 72 717
rect 85 669 101 717
rect 168 669 184 717
rect 195 669 211 717
rect 258 669 274 717
rect 285 669 301 717
rect 313 669 329 717
rect 340 669 356 717
rect 56 565 72 613
rect 85 565 101 613
rect 113 565 129 613
rect 166 565 182 613
rect 202 565 218 613
rect 258 565 274 613
rect 285 565 301 613
rect 56 487 72 535
rect 85 487 101 535
rect 56 408 72 456
rect 85 408 101 456
rect 168 487 184 535
rect 195 487 211 535
rect 258 487 274 535
rect 285 487 301 535
rect 168 408 184 456
rect 195 408 211 456
rect 250 408 266 456
rect 477 669 493 717
rect 504 669 520 717
rect 347 565 363 613
rect 403 565 419 613
rect 431 565 447 613
rect 460 565 476 613
rect 345 454 361 502
rect 378 454 394 502
rect 460 454 476 502
<< psubstratetap >>
rect 10 67 26 83
rect 38 67 54 83
rect 66 67 82 83
rect 94 67 110 83
rect 122 67 138 83
rect 150 67 166 83
rect 178 67 194 83
rect 206 67 222 83
rect 234 67 250 83
rect 262 67 278 83
rect 290 67 306 83
rect 318 67 334 83
rect 346 67 362 83
rect 374 67 390 83
rect 402 67 418 83
rect 430 67 446 83
rect 458 67 474 83
rect 486 67 502 83
<< nsubstratetap >>
rect 13 736 29 752
rect 41 736 57 752
rect 69 736 85 752
rect 97 736 113 752
rect 125 736 141 752
rect 153 736 169 752
rect 181 736 197 752
rect 209 736 225 752
rect 237 736 253 752
rect 265 736 281 752
rect 293 736 309 752
rect 321 736 337 752
rect 349 736 365 752
rect 377 736 393 752
rect 405 736 421 752
rect 433 736 449 752
rect 461 736 477 752
rect 489 736 505 752
<< metal1 >>
rect 0 782 528 792
rect 0 762 528 772
rect 0 736 13 752
rect 29 736 41 752
rect 57 736 69 752
rect 85 736 97 752
rect 113 736 125 752
rect 141 736 153 752
rect 169 736 181 752
rect 197 736 209 752
rect 225 736 237 752
rect 253 736 265 752
rect 281 736 293 752
rect 309 736 321 752
rect 337 736 349 752
rect 365 736 377 752
rect 393 736 405 752
rect 421 736 433 752
rect 449 736 461 752
rect 477 736 489 752
rect 505 736 528 752
rect 0 727 528 736
rect 6 555 16 727
rect 59 717 69 727
rect 316 717 326 727
rect 507 717 517 727
rect 101 688 168 698
rect 211 688 258 698
rect 356 688 390 698
rect 406 688 453 698
rect 467 688 477 698
rect 29 656 39 669
rect 29 646 65 656
rect 91 649 278 659
rect 91 613 101 649
rect 116 626 182 636
rect 116 613 126 626
rect 208 613 218 649
rect 268 633 278 649
rect 288 656 298 669
rect 288 646 326 656
rect 445 649 486 659
rect 268 623 363 633
rect 406 623 446 633
rect 288 613 298 623
rect 406 613 416 623
rect 476 603 486 649
rect 59 555 69 565
rect 116 555 126 565
rect 169 555 179 565
rect 260 555 270 565
rect 347 555 357 565
rect 6 545 357 555
rect 59 535 69 545
rect 260 535 270 545
rect 101 506 168 516
rect 211 506 238 516
rect 59 477 69 487
rect 228 477 238 506
rect 347 522 357 545
rect 431 522 441 565
rect 301 506 333 516
rect 347 512 441 522
rect 323 483 333 506
rect 381 502 391 512
rect 59 467 208 477
rect 228 467 312 477
rect 323 473 345 483
rect 59 456 69 467
rect 198 456 208 467
rect 101 427 168 437
rect 148 398 158 427
rect 266 427 276 437
rect 302 418 312 467
rect 476 473 486 483
rect 348 444 358 454
rect 348 434 446 444
rect 302 408 358 418
rect 148 388 418 398
rect 198 368 208 388
rect 99 344 168 354
rect 302 368 358 378
rect 59 328 69 338
rect 59 318 223 328
rect 266 328 276 338
rect 59 288 69 318
rect 302 308 312 368
rect 384 361 446 371
rect 384 331 394 361
rect 409 341 486 351
rect 409 331 419 341
rect 463 331 473 341
rect 123 298 312 308
rect 323 311 345 321
rect 123 278 133 298
rect 99 268 168 278
rect 323 278 333 311
rect 436 291 446 301
rect 301 268 333 278
rect 347 281 446 291
rect 59 248 69 258
rect 198 248 208 258
rect 261 248 271 258
rect 347 248 357 281
rect 6 238 357 248
rect 421 238 431 281
rect 6 92 16 238
rect 59 228 69 238
rect 99 208 168 218
rect 211 208 258 218
rect 301 208 321 218
rect 311 198 321 208
rect 384 198 394 208
rect 311 188 358 198
rect 91 178 298 188
rect 384 188 446 198
rect 29 155 65 165
rect 29 132 39 155
rect 91 132 101 178
rect 143 155 181 165
rect 143 132 153 155
rect 208 132 218 178
rect 288 168 326 178
rect 288 132 298 168
rect 316 142 390 152
rect 316 132 326 142
rect 476 166 486 218
rect 442 156 486 166
rect 356 112 453 122
rect 467 112 477 122
rect 56 92 66 102
rect 116 92 126 102
rect 171 92 181 102
rect 261 92 271 102
rect 507 92 517 102
rect 0 83 528 92
rect 0 67 10 83
rect 26 67 38 83
rect 54 67 66 83
rect 82 67 94 83
rect 110 67 122 83
rect 138 67 150 83
rect 166 67 178 83
rect 194 67 206 83
rect 222 67 234 83
rect 250 67 262 83
rect 278 67 290 83
rect 306 67 318 83
rect 334 67 346 83
rect 362 67 374 83
rect 390 67 402 83
rect 418 67 430 83
rect 446 67 458 83
rect 474 67 486 83
rect 502 67 528 83
rect 0 47 528 57
rect 0 27 528 37
rect 0 7 528 17
<< m2contact >>
rect 453 685 467 700
rect 431 649 445 663
rect 367 541 381 555
rect 392 541 406 555
rect 451 541 465 555
rect 43 384 57 398
rect 128 364 142 378
rect 237 364 251 378
rect 367 248 381 262
rect 392 248 406 262
rect 451 248 465 262
rect 428 154 442 168
rect 453 110 467 124
<< metal2 >>
rect 48 398 60 799
rect 57 384 60 398
rect 48 0 60 384
rect 120 378 132 799
rect 240 378 252 799
rect 432 722 444 799
rect 430 710 444 722
rect 430 663 442 710
rect 456 700 468 799
rect 467 697 468 700
rect 467 685 514 697
rect 430 661 431 663
rect 120 364 128 378
rect 251 364 252 378
rect 120 0 132 364
rect 240 0 252 364
rect 343 649 431 661
rect 343 168 355 649
rect 368 262 380 541
rect 393 262 405 541
rect 452 262 464 541
rect 343 156 428 168
rect 429 100 441 154
rect 467 122 468 124
rect 502 122 514 685
rect 467 110 514 122
rect 429 88 444 100
rect 432 0 444 88
rect 456 0 468 110
<< labels >>
rlabel metal2 48 0 60 0 1 A
rlabel metal2 120 0 132 0 1 B
rlabel metal2 240 0 252 0 1 Cin
rlabel metal2 432 0 444 0 1 S
rlabel metal2 456 0 468 0 1 Cout
rlabel metal2 48 799 60 799 5 A
rlabel metal2 456 799 468 799 5 Cout
rlabel metal2 432 799 444 799 5 S
rlabel metal2 240 799 252 799 5 Cin
rlabel metal2 120 799 132 799 5 B
rlabel metal1 528 27 528 37 7 Test
rlabel metal1 528 47 528 57 7 Clock
rlabel metal1 528 67 528 92 7 GND!
rlabel metal1 0 27 0 37 3 Test
rlabel metal1 0 47 0 57 3 Clock
rlabel metal1 0 67 0 92 3 GND!
rlabel metal1 528 727 528 752 7 Vdd!
rlabel metal1 528 782 528 792 7 ScanReturn
rlabel metal1 0 727 0 752 3 Vdd!
rlabel metal1 0 782 0 792 3 ScanReturn
rlabel metal1 0 762 0 772 3 Scan
rlabel metal1 528 762 528 772 7 Scan
rlabel metal1 0 7 0 17 3 nReset
rlabel metal1 528 7 528 17 7 nReset
<< end >>
