magic
tech c035u
timestamp 1385928057
<< nwell >>
rect 0 402 80 746
<< polysilicon >>
rect 60 756 62 772
rect 55 480 62 756
rect 55 362 62 432
rect 55 324 62 332
<< ndiffusion >>
rect 53 332 55 362
rect 62 332 64 362
<< pdiffusion >>
rect 53 432 55 480
rect 62 432 64 480
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 92 86
<< nohmic >>
rect 0 736 6 746
rect 22 736 34 746
<< ntransistor >>
rect 55 332 62 362
<< ptransistor >>
rect 55 432 62 480
<< polycontact >>
rect 44 756 60 772
<< ndiffcontact >>
rect 37 332 53 362
rect 64 332 80 362
<< pdiffcontact >>
rect 37 432 53 480
rect 64 432 80 480
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
<< nsubstratetap >>
rect 6 730 22 746
rect 34 730 50 746
<< metal1 >>
rect 0 782 80 792
rect 0 759 44 769
rect 0 730 6 746
rect 22 730 34 746
rect 50 730 53 746
rect 0 721 53 730
rect 37 480 53 721
rect 70 480 80 782
rect 70 362 80 432
rect 37 101 53 332
rect 0 92 92 101
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 92 92
<< m2contact >>
rect 92 76 292 101
<< metal2 >>
rect 92 101 292 799
rect 92 0 292 76
<< labels >>
rlabel metal2 92 799 292 799 5 GND!
rlabel metal2 92 0 292 0 1 GND!
rlabel metal1 0 759 0 769 7 Scan
rlabel metal1 0 721 0 746 3 Vdd!
rlabel metal1 0 782 0 792 3 nScan
rlabel metal1 0 76 0 101 7 GND!
<< end >>
