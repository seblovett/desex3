magic
tech c035u
timestamp 1385031005
<< nwell >>
rect 0 481 288 780
<< polysilicon >>
rect 216 669 221 685
rect 28 659 35 667
rect 58 659 65 667
rect 88 659 95 667
rect 132 659 139 667
rect 162 659 169 667
rect 189 659 196 667
rect 216 659 223 669
rect 28 372 35 611
rect 58 541 65 611
rect 88 527 95 611
rect 132 541 139 611
rect 88 511 93 527
rect 58 378 65 493
rect 28 236 35 356
rect 58 332 65 362
rect 88 332 95 511
rect 132 378 139 493
rect 162 378 169 611
rect 189 489 196 611
rect 132 332 139 362
rect 88 316 93 332
rect 58 236 65 306
rect 88 236 95 316
rect 132 236 139 306
rect 162 236 169 362
rect 189 352 196 473
rect 189 236 196 336
rect 216 236 223 611
rect 246 571 251 587
rect 246 541 253 571
rect 246 332 253 493
rect 246 276 253 306
rect 251 260 253 276
rect 28 202 35 210
rect 58 202 65 210
rect 88 202 95 210
rect 132 202 139 210
rect 162 202 169 210
rect 189 202 196 210
rect 216 202 223 210
<< ndiffusion >>
rect 56 306 58 332
rect 65 306 67 332
rect 130 306 132 332
rect 139 306 141 332
rect 244 306 246 332
rect 253 306 255 332
rect 26 210 28 236
rect 35 210 58 236
rect 65 210 67 236
rect 83 210 88 236
rect 95 210 114 236
rect 130 210 132 236
rect 139 210 162 236
rect 169 210 171 236
rect 187 210 189 236
rect 196 210 216 236
rect 223 210 225 236
<< pdiffusion >>
rect 26 611 28 659
rect 35 611 40 659
rect 56 611 58 659
rect 65 611 67 659
rect 83 611 88 659
rect 95 611 114 659
rect 130 611 132 659
rect 139 611 141 659
rect 157 611 162 659
rect 169 611 171 659
rect 187 611 189 659
rect 196 611 198 659
rect 214 611 216 659
rect 223 611 225 659
rect 56 493 58 541
rect 65 493 67 541
rect 130 493 132 541
rect 139 493 141 541
rect 244 493 246 541
rect 253 493 255 541
<< pohmic >>
rect 0 76 6 86
rect 22 76 34 86
rect 50 76 62 86
rect 78 76 90 86
rect 106 76 118 86
rect 134 76 146 86
rect 162 76 174 86
rect 190 76 202 86
rect 218 76 230 86
rect 246 76 258 86
rect 274 76 288 86
rect 0 73 288 76
<< nohmic >>
rect 0 731 288 734
rect 0 724 6 731
rect 22 724 34 731
rect 50 724 62 731
rect 78 724 90 731
rect 106 724 118 731
rect 134 724 146 731
rect 162 724 174 731
rect 190 724 202 731
rect 218 724 230 731
rect 246 724 258 731
rect 274 724 288 731
<< ntransistor >>
rect 58 306 65 332
rect 132 306 139 332
rect 246 306 253 332
rect 28 210 35 236
rect 58 210 65 236
rect 88 210 95 236
rect 132 210 139 236
rect 162 210 169 236
rect 189 210 196 236
rect 216 210 223 236
<< ptransistor >>
rect 28 611 35 659
rect 58 611 65 659
rect 88 611 95 659
rect 132 611 139 659
rect 162 611 169 659
rect 189 611 196 659
rect 216 611 223 659
rect 58 493 65 541
rect 132 493 139 541
rect 246 493 253 541
<< polycontact >>
rect 221 669 237 685
rect 93 511 109 527
rect 24 356 40 372
rect 54 362 70 378
rect 180 473 196 489
rect 127 362 143 378
rect 158 362 174 378
rect 93 316 109 332
rect 180 336 196 352
rect 251 571 267 587
rect 235 260 251 276
<< ndiffcontact >>
rect 40 306 56 332
rect 67 306 83 332
rect 114 306 130 332
rect 141 306 157 332
rect 228 306 244 332
rect 255 306 271 332
rect 10 210 26 236
rect 67 210 83 236
rect 114 210 130 236
rect 171 210 187 236
rect 225 210 241 236
<< pdiffcontact >>
rect 9 611 26 659
rect 40 611 56 659
rect 67 611 83 659
rect 114 611 130 659
rect 141 611 157 659
rect 171 611 187 659
rect 198 611 214 659
rect 225 611 241 659
rect 40 493 56 541
rect 67 493 83 541
rect 114 493 130 541
rect 141 493 157 541
rect 228 493 244 541
rect 255 493 271 541
<< psubstratetap >>
rect 6 76 22 92
rect 34 76 50 92
rect 62 76 78 92
rect 90 76 106 92
rect 118 76 134 92
rect 146 76 162 92
rect 174 76 190 92
rect 202 76 218 92
rect 230 76 246 92
rect 258 76 274 92
<< nsubstratetap >>
rect 6 715 22 731
rect 34 715 50 731
rect 62 715 78 731
rect 90 715 106 731
rect 118 715 134 731
rect 146 715 162 731
rect 174 715 190 731
rect 202 715 218 731
rect 230 715 246 731
rect 258 715 274 731
<< metal1 >>
rect 0 770 288 780
rect 0 747 174 757
rect 252 747 288 757
rect 0 731 288 734
rect 0 715 6 731
rect 22 715 34 731
rect 50 715 62 731
rect 78 715 90 731
rect 106 715 118 731
rect 134 715 146 731
rect 162 715 174 731
rect 190 715 202 731
rect 218 715 230 731
rect 246 715 258 731
rect 274 715 288 731
rect 0 709 288 715
rect 9 659 26 709
rect 67 659 83 709
rect 93 689 211 699
rect 15 561 26 611
rect 43 601 53 611
rect 93 601 103 689
rect 120 669 184 679
rect 120 659 130 669
rect 174 659 184 669
rect 201 659 211 689
rect 43 591 103 601
rect 144 581 154 611
rect 174 601 184 611
rect 228 601 238 611
rect 174 591 238 601
rect 144 571 251 581
rect 15 551 238 561
rect 40 541 50 551
rect 145 541 157 551
rect 109 511 114 527
rect 228 541 238 551
rect 73 483 83 493
rect 73 473 180 483
rect 261 385 271 493
rect 70 364 72 378
rect 120 362 127 376
rect 261 375 288 385
rect 73 342 180 352
rect 73 332 83 342
rect 261 332 271 375
rect 109 316 114 332
rect 46 296 56 306
rect 147 296 157 306
rect 228 296 238 306
rect 46 286 271 296
rect 13 266 235 276
rect 13 236 23 266
rect 70 246 150 256
rect 70 236 80 246
rect 114 98 130 210
rect 140 200 150 246
rect 174 236 184 266
rect 228 200 238 210
rect 140 190 238 200
rect 261 98 271 286
rect 0 92 288 98
rect 0 76 6 92
rect 22 76 34 92
rect 50 76 62 92
rect 78 76 90 92
rect 106 76 118 92
rect 134 76 146 92
rect 162 76 174 92
rect 190 76 202 92
rect 218 76 230 92
rect 246 76 258 92
rect 274 76 288 92
rect 0 73 288 76
rect 0 50 288 60
rect 0 27 106 37
rect 120 27 288 37
rect 0 4 288 14
<< m2contact >>
rect 174 745 188 759
rect 238 746 252 760
rect 237 671 251 685
rect 72 364 87 378
rect 106 362 120 376
rect 174 364 188 378
rect 24 342 38 356
rect 106 25 120 39
<< metal2 >>
rect 24 356 36 783
rect 75 378 87 783
rect 175 731 187 745
rect 174 715 187 731
rect 175 378 187 715
rect 239 685 251 746
rect 24 0 36 342
rect 75 0 87 364
rect 107 39 119 362
<< labels >>
rlabel metal1 0 73 0 98 3 GND!
rlabel metal1 0 27 0 37 3 Test
rlabel metal1 0 4 0 14 2 nReset
rlabel metal1 0 50 0 60 3 Clock
rlabel metal2 24 0 36 0 1 D
rlabel metal2 75 0 87 0 1 Load
rlabel metal1 288 50 288 60 7 Clock
rlabel metal1 288 27 288 37 7 Test
rlabel metal1 288 4 288 14 8 nReset
rlabel metal1 288 73 288 98 7 GND!
rlabel metal1 0 770 0 780 3 ScanReturn
rlabel metal1 0 747 0 757 3 SDI
rlabel metal1 0 709 0 734 3 Vdd!
rlabel metal1 288 709 288 734 1 Vdd!
rlabel metal1 288 747 288 757 7 Q
rlabel metal1 288 770 288 780 7 ScanReturn
rlabel metal2 24 783 36 783 5 D
rlabel metal2 75 783 87 783 5 Load
rlabel metal1 288 375 288 385 7 M
<< end >>
