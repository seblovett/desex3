magic
tech c035u
timestamp 1384897405
<< nwell >>
rect 1929 290 2079 502
<< metal1 >>
rect 1929 540 2079 550
rect 3519 540 3545 550
rect 1929 516 2079 526
rect 1929 477 2079 502
rect 1929 162 2079 187
rect 3519 162 3545 187
rect 1929 138 1976 148
rect 1990 138 2079 148
rect 1929 114 2014 124
rect 2028 114 2079 124
rect 1929 90 2055 100
rect 2069 90 2079 100
rect 2070 66 2462 76
rect 2476 66 2582 76
rect 2596 66 2702 76
rect 2029 44 2822 54
rect 2836 44 2942 54
rect 2956 44 3062 54
rect 1991 22 2101 32
rect 2115 22 2222 32
rect 2236 22 2342 32
<< m2contact >>
rect 1976 136 1990 150
rect 2014 112 2028 126
rect 2055 88 2069 102
rect 2056 64 2070 78
rect 2462 64 2476 78
rect 2582 64 2596 78
rect 2702 65 2716 79
rect 2015 44 2029 58
rect 2822 42 2836 56
rect 2942 43 2956 57
rect 3062 41 3076 55
rect 1977 20 1991 34
rect 2101 20 2115 34
rect 2222 20 2236 34
rect 2342 20 2356 34
<< metal2 >>
rect 0 586 200 653
rect 223 622 235 653
rect 223 610 3435 622
rect 223 586 235 610
rect 3183 554 3195 610
rect 3303 554 3315 610
rect 3423 554 3435 610
rect 0 0 200 77
rect 223 0 235 77
rect 247 0 259 77
rect 271 0 283 77
rect 295 0 307 77
rect 1978 34 1990 136
rect 2016 58 2028 112
rect 2056 78 2069 88
rect 1978 0 1990 20
rect 2016 0 2028 44
rect 2057 0 2069 64
rect 2103 34 2115 89
rect 2223 34 2235 89
rect 2343 34 2355 89
rect 2463 78 2475 89
rect 2583 78 2595 89
rect 2703 79 2715 89
rect 2823 56 2835 89
rect 2943 57 2955 89
rect 3063 55 3075 89
use leftbuf leftbuf_0
timestamp 1384893035
transform 1 0 0 0 1 77
box 0 0 1929 509
use inv inv_0
timestamp 1384893302
transform 1 0 2079 0 1 89
box 0 0 120 465
use inv inv_1
timestamp 1384893302
transform 1 0 2199 0 1 89
box 0 0 120 465
use inv inv_2
timestamp 1384893302
transform 1 0 2319 0 1 89
box 0 0 120 465
use inv inv_3
timestamp 1384893302
transform 1 0 2439 0 1 89
box 0 0 120 465
use inv inv_4
timestamp 1384893302
transform 1 0 2559 0 1 89
box 0 0 120 465
use inv inv_5
timestamp 1384893302
transform 1 0 2679 0 1 89
box 0 0 120 465
use inv inv_6
timestamp 1384893302
transform 1 0 2799 0 1 89
box 0 0 120 465
use inv inv_7
timestamp 1384893302
transform 1 0 2919 0 1 89
box 0 0 120 465
use inv inv_8
timestamp 1384893302
transform 1 0 3039 0 1 89
box 0 0 120 465
use inv inv_9
timestamp 1384893302
transform 1 0 3159 0 1 89
box 0 0 120 465
use inv inv_10
timestamp 1384893302
transform 1 0 3279 0 1 89
box 0 0 120 465
use inv inv_11
timestamp 1384893302
transform 1 0 3399 0 1 89
box 0 0 120 465
<< labels >>
rlabel metal2 1978 0 1990 0 1 ClockOut
rlabel metal2 2016 0 2028 0 1 TestOut
rlabel metal2 2057 0 2069 0 1 ResetOut
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 247 0 259 0 1 Test
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 295 0 307 0 1 nReset
rlabel metal2 223 653 235 653 5 SDO
rlabel metal2 0 653 200 653 5 Vdd!
rlabel metal1 3545 162 3545 187 7 GND!
rlabel metal1 3545 540 3545 550 7 nSDO
rlabel metal2 0 0 200 0 1 Vdd!
<< end >>
