magic
tech c035u
timestamp 1386006472
<< nwell >>
rect 202 402 1464 746
rect 405 401 451 402
rect 742 401 788 402
rect 1079 401 1125 402
<< polysilicon >>
rect 538 692 545 700
rect 565 692 572 700
rect 592 692 599 700
rect 619 692 626 700
rect 875 692 882 700
rect 902 692 909 700
rect 929 692 936 700
rect 956 692 963 700
rect 1212 692 1219 700
rect 1239 692 1246 700
rect 1266 692 1273 700
rect 1293 692 1300 700
rect 480 614 487 622
rect 507 614 514 622
rect 425 559 432 567
rect 370 460 377 468
rect 817 614 824 622
rect 844 614 851 622
rect 762 559 769 567
rect 707 460 714 468
rect 1154 614 1161 622
rect 1181 614 1188 622
rect 1099 559 1106 567
rect 1044 460 1051 468
rect 1394 516 1396 532
rect 1389 471 1396 516
rect 370 388 377 402
rect 425 388 432 402
rect 480 389 487 402
rect 375 372 377 388
rect 430 372 432 388
rect 485 385 487 389
rect 507 385 514 402
rect 538 389 545 402
rect 485 378 514 385
rect 485 373 487 378
rect 543 385 545 389
rect 565 385 572 402
rect 592 385 599 402
rect 619 385 626 402
rect 707 388 714 402
rect 762 388 769 402
rect 817 389 824 402
rect 543 378 626 385
rect 543 373 545 378
rect 370 362 377 372
rect 425 362 432 372
rect 480 362 487 373
rect 538 362 545 373
rect 565 362 572 378
rect 712 372 714 388
rect 767 372 769 388
rect 822 385 824 389
rect 844 385 851 402
rect 875 389 882 402
rect 822 378 851 385
rect 822 373 824 378
rect 880 385 882 389
rect 902 385 909 402
rect 929 385 936 402
rect 956 385 963 402
rect 1044 388 1051 402
rect 1099 388 1106 402
rect 1154 389 1161 402
rect 880 378 963 385
rect 880 373 882 378
rect 707 362 714 372
rect 762 362 769 372
rect 817 362 824 373
rect 875 362 882 373
rect 902 362 909 378
rect 1049 372 1051 388
rect 1104 372 1106 388
rect 1159 385 1161 389
rect 1181 385 1188 402
rect 1212 389 1219 402
rect 1159 378 1188 385
rect 1159 373 1161 378
rect 1217 385 1219 389
rect 1239 385 1246 402
rect 1266 385 1273 402
rect 1293 385 1300 402
rect 1217 378 1300 385
rect 1217 373 1219 378
rect 1044 362 1051 372
rect 1099 362 1106 372
rect 1154 362 1161 373
rect 1212 362 1219 373
rect 1239 362 1246 378
rect 1389 377 1396 423
rect 370 334 377 342
rect 425 300 432 308
rect 480 208 487 216
rect 707 334 714 342
rect 762 300 769 308
rect 817 208 824 216
rect 1044 334 1051 342
rect 1099 300 1106 308
rect 1154 208 1161 216
rect 1389 339 1396 347
rect 538 154 545 162
rect 565 154 572 162
rect 875 154 882 162
rect 902 154 909 162
rect 1212 154 1219 162
rect 1239 154 1246 162
<< ndiffusion >>
rect 368 342 370 362
rect 377 342 379 362
rect 423 308 425 362
rect 432 308 434 362
rect 478 216 480 362
rect 487 216 489 362
rect 536 162 538 362
rect 545 162 547 362
rect 563 162 565 362
rect 572 162 574 362
rect 705 342 707 362
rect 714 342 716 362
rect 760 308 762 362
rect 769 308 771 362
rect 815 216 817 362
rect 824 216 826 362
rect 873 162 875 362
rect 882 162 884 362
rect 900 162 902 362
rect 909 162 911 362
rect 1042 342 1044 362
rect 1051 342 1053 362
rect 1097 308 1099 362
rect 1106 308 1108 362
rect 1152 216 1154 362
rect 1161 216 1163 362
rect 1210 162 1212 362
rect 1219 162 1221 362
rect 1237 162 1239 362
rect 1246 162 1248 362
rect 1387 347 1389 377
rect 1396 347 1398 377
<< pdiffusion >>
rect 368 402 370 460
rect 377 402 379 460
rect 423 402 425 559
rect 432 402 434 559
rect 478 402 480 614
rect 487 402 489 614
rect 505 402 507 614
rect 514 402 516 614
rect 536 402 538 692
rect 545 402 547 692
rect 563 402 565 692
rect 572 402 574 692
rect 590 402 592 692
rect 599 402 601 692
rect 617 402 619 692
rect 626 402 628 692
rect 705 402 707 460
rect 714 402 716 460
rect 760 402 762 559
rect 769 402 771 559
rect 815 402 817 614
rect 824 402 826 614
rect 842 402 844 614
rect 851 402 853 614
rect 873 402 875 692
rect 882 402 884 692
rect 900 402 902 692
rect 909 402 911 692
rect 927 402 929 692
rect 936 402 938 692
rect 954 402 956 692
rect 963 402 965 692
rect 1042 402 1044 460
rect 1051 402 1053 460
rect 1097 402 1099 559
rect 1106 402 1108 559
rect 1152 402 1154 614
rect 1161 402 1163 614
rect 1179 402 1181 614
rect 1188 402 1190 614
rect 1210 402 1212 692
rect 1219 402 1221 692
rect 1237 402 1239 692
rect 1246 402 1248 692
rect 1264 402 1266 692
rect 1273 402 1275 692
rect 1291 402 1293 692
rect 1300 402 1302 692
rect 1387 423 1389 471
rect 1396 423 1398 471
<< pohmic >>
rect 320 76 326 86
rect 342 76 354 86
rect 370 76 382 86
rect 398 76 410 86
rect 426 76 438 86
rect 454 76 466 86
rect 482 76 494 86
rect 510 76 522 86
rect 538 76 550 86
rect 567 76 579 86
rect 595 76 607 86
rect 623 76 635 86
rect 651 76 663 86
rect 679 76 691 86
rect 707 76 719 86
rect 735 76 747 86
rect 763 76 775 86
rect 791 76 803 86
rect 819 76 831 86
rect 847 76 859 86
rect 875 76 887 86
rect 904 76 916 86
rect 932 76 944 86
rect 960 76 972 86
rect 988 76 1000 86
rect 1016 76 1028 86
rect 1044 76 1056 86
rect 1072 76 1084 86
rect 1100 76 1112 86
rect 1128 76 1140 86
rect 1156 76 1168 86
rect 1184 76 1196 86
rect 1212 76 1224 86
rect 1241 76 1253 86
rect 1269 76 1281 86
rect 1297 76 1309 86
rect 1325 76 1337 86
rect 1353 76 1365 86
rect 1381 76 1393 86
rect 1409 76 1421 86
rect 1437 76 1464 86
<< nohmic >>
rect 202 736 214 746
rect 230 736 242 746
rect 258 736 270 746
rect 286 736 298 746
rect 314 736 326 746
rect 342 736 354 746
rect 370 736 382 746
rect 398 736 410 746
rect 426 736 438 746
rect 454 736 466 746
rect 482 736 494 746
rect 510 736 522 746
rect 538 736 550 746
rect 567 736 579 746
rect 595 736 607 746
rect 623 736 635 746
rect 651 736 663 746
rect 679 736 691 746
rect 707 736 719 746
rect 735 736 747 746
rect 763 736 775 746
rect 791 736 803 746
rect 819 736 831 746
rect 847 736 859 746
rect 875 736 887 746
rect 904 736 916 746
rect 932 736 944 746
rect 960 736 972 746
rect 988 736 1000 746
rect 1016 736 1028 746
rect 1044 736 1056 746
rect 1072 736 1084 746
rect 1100 736 1112 746
rect 1128 736 1140 746
rect 1156 736 1168 746
rect 1184 736 1196 746
rect 1212 736 1224 746
rect 1241 736 1253 746
rect 1269 736 1281 746
rect 1297 736 1309 746
rect 1325 736 1337 746
rect 1353 736 1365 746
rect 1381 736 1393 746
rect 1409 736 1421 746
rect 1437 736 1464 746
<< ntransistor >>
rect 370 342 377 362
rect 425 308 432 362
rect 480 216 487 362
rect 538 162 545 362
rect 565 162 572 362
rect 707 342 714 362
rect 762 308 769 362
rect 817 216 824 362
rect 875 162 882 362
rect 902 162 909 362
rect 1044 342 1051 362
rect 1099 308 1106 362
rect 1154 216 1161 362
rect 1212 162 1219 362
rect 1239 162 1246 362
rect 1389 347 1396 377
<< ptransistor >>
rect 370 402 377 460
rect 425 402 432 559
rect 480 402 487 614
rect 507 402 514 614
rect 538 402 545 692
rect 565 402 572 692
rect 592 402 599 692
rect 619 402 626 692
rect 707 402 714 460
rect 762 402 769 559
rect 817 402 824 614
rect 844 402 851 614
rect 875 402 882 692
rect 902 402 909 692
rect 929 402 936 692
rect 956 402 963 692
rect 1044 402 1051 460
rect 1099 402 1106 559
rect 1154 402 1161 614
rect 1181 402 1188 614
rect 1212 402 1219 692
rect 1239 402 1246 692
rect 1266 402 1273 692
rect 1293 402 1300 692
rect 1389 423 1396 471
<< polycontact >>
rect 1378 516 1394 532
rect 359 372 375 388
rect 414 372 430 388
rect 469 373 485 389
rect 527 373 543 389
rect 696 372 712 388
rect 751 372 767 388
rect 806 373 822 389
rect 864 373 880 389
rect 1033 372 1049 388
rect 1088 372 1104 388
rect 1143 373 1159 389
rect 1201 373 1217 389
<< ndiffcontact >>
rect 352 342 368 362
rect 379 342 395 362
rect 407 308 423 362
rect 434 308 450 362
rect 462 216 478 362
rect 489 216 505 362
rect 520 162 536 362
rect 547 162 563 362
rect 574 162 590 362
rect 689 342 705 362
rect 716 342 732 362
rect 744 308 760 362
rect 771 308 787 362
rect 799 216 815 362
rect 826 216 842 362
rect 857 162 873 362
rect 884 162 900 362
rect 911 162 927 362
rect 1026 342 1042 362
rect 1053 342 1069 362
rect 1081 308 1097 362
rect 1108 308 1124 362
rect 1136 216 1152 362
rect 1163 216 1179 362
rect 1194 162 1210 362
rect 1221 162 1237 362
rect 1248 162 1264 362
rect 1371 347 1387 377
rect 1398 347 1414 377
<< pdiffcontact >>
rect 519 614 536 692
rect 352 402 368 460
rect 379 402 395 460
rect 407 402 423 559
rect 434 402 450 559
rect 462 402 478 614
rect 489 402 505 614
rect 516 402 536 614
rect 547 402 563 692
rect 574 402 590 692
rect 601 402 617 692
rect 628 402 644 692
rect 856 614 873 692
rect 689 402 705 460
rect 716 402 732 460
rect 744 402 760 559
rect 771 402 787 559
rect 799 402 815 614
rect 826 402 842 614
rect 853 402 873 614
rect 884 402 900 692
rect 911 402 927 692
rect 938 402 954 692
rect 965 402 981 692
rect 1193 614 1210 692
rect 1026 402 1042 460
rect 1053 402 1069 460
rect 1081 402 1097 559
rect 1108 402 1124 559
rect 1136 402 1152 614
rect 1163 402 1179 614
rect 1190 402 1210 614
rect 1221 402 1237 692
rect 1248 402 1264 692
rect 1275 402 1291 692
rect 1302 402 1318 692
rect 1371 423 1387 471
rect 1398 423 1414 471
<< psubstratetap >>
rect 326 76 342 92
rect 354 76 370 92
rect 382 76 398 92
rect 410 76 426 92
rect 438 76 454 92
rect 466 76 482 92
rect 494 76 510 92
rect 522 76 538 92
rect 550 76 567 92
rect 579 76 595 92
rect 607 76 623 92
rect 635 76 651 92
rect 663 76 679 92
rect 691 76 707 92
rect 719 76 735 92
rect 747 76 763 92
rect 775 76 791 92
rect 803 76 819 92
rect 831 76 847 92
rect 859 76 875 92
rect 887 76 904 92
rect 916 76 932 92
rect 944 76 960 92
rect 972 76 988 92
rect 1000 76 1016 92
rect 1028 76 1044 92
rect 1056 76 1072 92
rect 1084 76 1100 92
rect 1112 76 1128 92
rect 1140 76 1156 92
rect 1168 76 1184 92
rect 1196 76 1212 92
rect 1224 76 1241 92
rect 1253 76 1269 92
rect 1281 76 1297 92
rect 1309 76 1325 92
rect 1337 76 1353 92
rect 1365 76 1381 92
rect 1393 76 1409 92
rect 1421 76 1437 92
<< nsubstratetap >>
rect 214 730 230 746
rect 242 730 258 746
rect 270 730 286 746
rect 298 730 314 746
rect 326 730 342 746
rect 354 730 370 746
rect 382 730 398 746
rect 410 730 426 746
rect 438 730 454 746
rect 466 730 482 746
rect 494 730 510 746
rect 522 730 538 746
rect 550 730 567 746
rect 579 730 595 746
rect 607 730 623 746
rect 635 730 651 746
rect 663 730 679 746
rect 691 730 707 746
rect 719 730 735 746
rect 747 730 763 746
rect 775 730 791 746
rect 803 730 819 746
rect 831 730 847 746
rect 859 730 875 746
rect 887 730 904 746
rect 916 730 932 746
rect 944 730 960 746
rect 972 730 988 746
rect 1000 730 1016 746
rect 1028 730 1044 746
rect 1056 730 1072 746
rect 1084 730 1100 746
rect 1112 730 1128 746
rect 1140 730 1156 746
rect 1168 730 1184 746
rect 1196 730 1212 746
rect 1224 730 1241 746
rect 1253 730 1269 746
rect 1281 730 1297 746
rect 1309 730 1325 746
rect 1337 730 1353 746
rect 1365 730 1381 746
rect 1393 730 1409 746
rect 1421 730 1437 746
<< metal1 >>
rect 185 756 200 792
rect 229 782 1356 792
rect 1400 782 1464 792
rect 229 759 1464 769
rect 200 730 214 746
rect 230 730 242 746
rect 258 730 270 746
rect 286 730 298 746
rect 314 730 326 746
rect 342 730 354 746
rect 370 730 382 746
rect 398 730 410 746
rect 426 730 438 746
rect 454 730 466 746
rect 482 730 494 746
rect 510 730 522 746
rect 538 730 550 746
rect 567 730 579 746
rect 595 730 607 746
rect 623 730 635 746
rect 651 730 663 746
rect 679 730 691 746
rect 707 730 719 746
rect 735 730 747 746
rect 763 730 775 746
rect 791 730 803 746
rect 819 730 831 746
rect 847 730 859 746
rect 875 730 887 746
rect 904 730 916 746
rect 932 730 944 746
rect 960 730 972 746
rect 988 730 1000 746
rect 1016 730 1028 746
rect 1044 730 1056 746
rect 1072 730 1084 746
rect 1100 730 1112 746
rect 1128 730 1140 746
rect 1156 730 1168 746
rect 1184 730 1196 746
rect 1212 730 1224 746
rect 1241 730 1253 746
rect 1269 730 1281 746
rect 1297 730 1309 746
rect 1325 730 1337 746
rect 1353 730 1365 746
rect 1381 730 1393 746
rect 1409 730 1421 746
rect 1437 730 1464 746
rect 200 721 1464 730
rect 352 460 368 721
rect 407 559 423 721
rect 462 614 478 721
rect 516 692 536 721
rect 574 692 590 721
rect 628 692 644 721
rect 516 614 519 692
rect 689 460 705 721
rect 744 559 760 721
rect 799 614 815 721
rect 853 692 873 721
rect 911 692 927 721
rect 965 692 981 721
rect 853 614 856 692
rect 1026 460 1042 721
rect 1081 559 1097 721
rect 1136 614 1152 721
rect 1190 692 1210 721
rect 1248 692 1264 721
rect 1302 692 1318 721
rect 1190 614 1193 692
rect 1380 532 1394 538
rect 1404 471 1414 721
rect 240 349 252 387
rect 277 375 359 385
rect 263 363 277 373
rect 385 385 395 402
rect 385 375 414 385
rect 385 362 395 375
rect 440 386 450 402
rect 440 376 469 386
rect 440 362 450 376
rect 495 386 505 402
rect 495 376 527 386
rect 495 362 505 376
rect 553 387 563 402
rect 607 389 617 402
rect 553 377 606 387
rect 553 362 563 377
rect 667 375 696 385
rect 722 385 732 402
rect 722 375 751 385
rect 722 362 732 375
rect 777 386 787 402
rect 777 376 806 386
rect 777 362 787 376
rect 832 386 842 402
rect 832 376 864 386
rect 832 362 842 376
rect 890 387 900 402
rect 944 389 954 402
rect 890 377 944 387
rect 890 362 900 377
rect 1022 375 1033 385
rect 1059 385 1069 402
rect 1059 375 1088 385
rect 1059 362 1069 375
rect 1114 386 1124 402
rect 1114 376 1143 386
rect 1114 362 1124 376
rect 1169 386 1179 402
rect 1169 376 1201 386
rect 1169 362 1179 376
rect 1227 387 1237 402
rect 1281 389 1291 402
rect 1227 377 1279 387
rect 1227 362 1237 377
rect 1371 377 1381 423
rect 352 101 368 342
rect 407 101 423 308
rect 462 101 478 216
rect 520 101 536 162
rect 574 101 590 162
rect 689 101 705 342
rect 744 101 760 308
rect 799 101 815 216
rect 857 101 873 162
rect 911 101 927 162
rect 1026 101 1042 342
rect 1081 101 1097 308
rect 1136 101 1152 216
rect 1194 101 1210 162
rect 1248 101 1264 162
rect 1398 101 1408 347
rect 320 92 1464 101
rect 320 76 326 92
rect 342 76 354 92
rect 370 76 382 92
rect 398 76 410 92
rect 426 76 438 92
rect 454 76 466 92
rect 482 76 494 92
rect 510 76 522 92
rect 538 76 550 92
rect 567 76 579 92
rect 595 76 607 92
rect 623 76 635 92
rect 651 76 663 92
rect 679 76 691 92
rect 707 76 719 92
rect 735 76 747 92
rect 763 76 775 92
rect 791 76 803 92
rect 819 76 831 92
rect 847 76 859 92
rect 875 76 887 92
rect 904 76 916 92
rect 932 76 944 92
rect 960 76 972 92
rect 988 76 1000 92
rect 1016 76 1028 92
rect 1044 76 1056 92
rect 1072 76 1084 92
rect 1100 76 1112 92
rect 1128 76 1140 92
rect 1156 76 1168 92
rect 1184 76 1196 92
rect 1212 76 1224 92
rect 1241 76 1253 92
rect 1269 76 1281 92
rect 1297 76 1309 92
rect 1325 76 1337 92
rect 1353 76 1365 92
rect 1381 76 1393 92
rect 1409 76 1421 92
rect 1437 76 1464 92
rect 216 4 228 67
rect 239 43 253 53
rect 620 53 1464 63
rect 253 30 653 40
rect 959 30 1464 40
rect 301 7 1009 17
rect 1033 7 1270 17
rect 1294 7 1304 17
rect 1318 7 1464 17
<< m2contact >>
rect 215 780 229 794
rect 1356 781 1370 795
rect 1386 781 1400 795
rect 215 756 229 770
rect 0 721 200 746
rect 1380 538 1394 552
rect 1357 457 1371 471
rect 263 373 277 387
rect 263 349 277 363
rect 606 375 620 389
rect 653 373 667 387
rect 944 375 958 389
rect 1008 373 1022 387
rect 1279 375 1293 389
rect 239 53 253 67
rect 606 51 620 65
rect 239 29 253 43
rect 653 28 667 42
rect 945 29 959 43
rect 239 5 253 19
rect 263 5 277 19
rect 287 5 301 19
rect 1009 5 1023 19
rect 1280 5 1294 19
rect 1304 5 1318 19
<< metal2 >>
rect 0 746 200 799
rect 216 794 228 799
rect 0 0 200 721
rect 216 0 228 756
rect 240 67 252 799
rect 264 387 276 799
rect 264 363 276 373
rect 240 43 252 53
rect 240 19 252 29
rect 264 19 276 349
rect 288 19 300 799
rect 1358 471 1370 781
rect 1386 552 1398 781
rect 1394 538 1398 552
rect 607 65 619 375
rect 654 42 666 373
rect 946 43 958 375
rect 1010 19 1022 373
rect 1281 19 1293 375
rect 1294 5 1304 19
rect 240 0 252 5
rect 264 0 276 5
rect 288 0 300 5
<< labels >>
rlabel metal2 0 799 200 799 5 Vdd!
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal1 1464 721 1464 746 7 Vdd!
rlabel metal1 1464 759 1464 769 7 SDI
rlabel metal1 1464 782 1464 792 7 nSDO
rlabel metal1 1464 53 1464 63 7 ClockOut
rlabel metal1 1464 30 1464 40 7 TestOut
rlabel metal1 1464 7 1464 17 7 nResetOut
rlabel metal1 1464 76 1464 101 7 GND!
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 288 799 300 799 5 nReset
rlabel metal2 240 799 252 799 5 Test
rlabel metal2 264 799 276 799 5 Clock
rlabel metal2 216 799 228 799 5 SDO
<< end >>
