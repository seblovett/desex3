magic
tech c035u
timestamp 1385631890
<< metal1 >>
rect 236 908 2660 918
rect 2674 908 2780 918
rect 2794 908 2900 918
rect 1443 865 1557 875
rect 2997 865 3077 875
rect 1443 842 1557 852
rect 2997 842 3077 852
rect 1443 804 1557 829
rect 2997 804 3077 829
rect 1443 159 1557 184
rect 2997 159 3077 184
rect 1443 136 1509 146
rect 1523 136 1557 146
rect 2997 136 3077 146
rect 1443 113 1486 123
rect 1500 113 1557 123
rect 2997 113 3077 123
rect 1443 90 1462 100
rect 1476 90 1557 100
rect 2997 90 3077 100
rect 1523 50 1580 60
rect 1594 50 1700 60
rect 1714 50 1820 60
rect 1500 28 1940 38
rect 1954 28 2060 38
rect 2074 28 2180 38
rect 1477 4 2300 14
rect 2314 4 2420 14
rect 2434 4 2540 14
<< m2contact >>
rect 222 907 236 921
rect 2660 906 2674 920
rect 2780 906 2794 920
rect 2900 906 2914 920
rect 1509 134 1523 148
rect 1486 110 1500 124
rect 1462 87 1476 101
rect 1509 50 1523 64
rect 1580 48 1594 62
rect 1700 48 1714 62
rect 1820 48 1834 62
rect 1486 26 1500 40
rect 1940 26 1954 40
rect 2060 26 2074 40
rect 2180 26 2194 40
rect 1463 2 1477 16
rect 2300 2 2314 16
rect 2420 2 2434 16
rect 2540 2 2554 16
<< metal2 >>
rect 223 921 235 934
rect 223 882 235 907
rect 2661 882 2673 906
rect 2781 882 2793 906
rect 2901 882 2913 906
rect 0 0 200 83
rect 223 0 235 83
rect 247 0 259 83
rect 271 0 283 83
rect 295 0 307 83
rect 1464 16 1476 87
rect 1487 40 1499 110
rect 1510 64 1522 134
rect 1581 62 1593 83
rect 1701 62 1713 83
rect 1821 62 1833 83
rect 1941 40 1953 83
rect 2061 40 2073 83
rect 2181 40 2193 83
rect 2301 16 2313 83
rect 2421 16 2433 83
rect 2541 16 2553 83
use leftbuf leftbuf_0
timestamp 1385631441
transform 1 0 0 0 1 93
box 0 -10 1443 789
use inv inv_0
timestamp 1385631115
transform 1 0 1557 0 1 83
box 0 0 120 799
use inv inv_1
timestamp 1385631115
transform 1 0 1677 0 1 83
box 0 0 120 799
use inv inv_2
timestamp 1385631115
transform 1 0 1797 0 1 83
box 0 0 120 799
use inv inv_3
timestamp 1385631115
transform 1 0 1917 0 1 83
box 0 0 120 799
use inv inv_4
timestamp 1385631115
transform 1 0 2037 0 1 83
box 0 0 120 799
use inv inv_5
timestamp 1385631115
transform 1 0 2157 0 1 83
box 0 0 120 799
use inv inv_6
timestamp 1385631115
transform 1 0 2277 0 1 83
box 0 0 120 799
use inv inv_7
timestamp 1385631115
transform 1 0 2397 0 1 83
box 0 0 120 799
use inv inv_8
timestamp 1385631115
transform 1 0 2517 0 1 83
box 0 0 120 799
use inv inv_9
timestamp 1385631115
transform 1 0 2637 0 1 83
box 0 0 120 799
use inv inv_10
timestamp 1385631115
transform 1 0 2757 0 1 83
box 0 0 120 799
use inv inv_11
timestamp 1385631115
transform 1 0 2877 0 1 83
box 0 0 120 799
<< labels >>
rlabel metal2 223 934 235 934 5 SDO
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 223 0 235 0 1 SDI
rlabel metal2 247 0 259 0 1 Test
rlabel metal2 271 0 283 0 1 Clock
rlabel metal2 295 0 307 0 1 nReset
rlabel metal1 3077 865 3077 875 7 nSDO
rlabel metal1 3077 842 3077 852 7 SDI
rlabel metal1 3077 804 3077 829 7 Vdd!
rlabel metal1 3077 90 3077 100 7 nResetOut
rlabel metal1 3077 113 3077 123 7 TestOut
rlabel metal1 3077 136 3077 146 7 ClockOut
rlabel metal1 3077 159 3077 184 7 GND!
<< end >>
